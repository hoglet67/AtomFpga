
package board_config_pack is

    constant G_CONFIG_DEBUGGER : boolean := true;

    constant G_CONFIG_VGA      : boolean := true;

end board_config_pack;


package body board_config_pack is

end board_config_pack;
