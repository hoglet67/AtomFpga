--
--Written by GowinSynthesis
--Product Version "V1.9.9 Beta"
--Thu May 11 17:52:08 2023

--Source file index table:
--file0 "\/disk1/home/dmb/gowin/v1.9.9beta/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\/disk1/home/dmb/gowin/v1.9.9beta/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
r9CEsN3Hgz//JHUvlMeZfgmQts6iFWnn7+wZf99REKtmm/5A/QEoed5v/lysn5s23E7x7vUZkZ3j
Z9uhVLk2kz5rxFYNPKyx8QD4UqK9ZebjMih8pHL9w55O0lHUaUXc9o/TCcLx/oIFy8gc26bHpbAo
2fmEbBmQ0UJuBk3DhcMT5XNYcL0M66x2k2yEXSm0hxqk4peLM/+3i7BjgzNKyBZCEGs+YHhHnDli
LzNOO47unlVoomOkIa3eADzM0w4G+QV40Rpo7/mF+oBfmT6veqUoP89m2WggXd0NMWKIGaD5N58P
GcYXF70hYZJN4Glup5h7mkj8H4nFCq8N0iSKmg==

`protect encoding=(enctype="base64", line_length=76, bytes=65280)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
qqJVEzFp6wSO+T1Baa3uT6w/s0ZqoS2heSOSam4mWy6msjtz3rznwU43tAdABZsVbH+9zCKg7O9i
/prhX+EdHO7gPZTIGuJRkVEGB4thKWxgaeIbV31NJFM/2VpCR3VjSU5SSlmQheqkcEoSmUvsMfUR
dECi3YE5rgeJKlGQHI76Uvv2fwIs52EN3cSysHOvjpIm4mLpiUAKr5ce1Wjs6YKqTKrEBWAa7QBf
QGU57EMXJIVFocPcd/4i1frbkvisMvuU5IFKLTYeBwYAaTEPHQl4ohSir+DjrfwRNpyUfVSR79XS
3yQ+UsU8Y55QSvbZ5fAfDcWXC/3FH+QkeXN6rJRDtSPJb3kZSply+3BsxNllKUSn3Tl3UUZr1GIT
AOmBCtyjejnW8xvAX8K/iYhRWuBJlT6PZLV3/0Hsdkb6tIWR+DAUa1qGlD3mqfek+VxN0GZyu6Vc
pyVy244uCmOMkIEUk1K/hMlt4XLhUj0f2WNHoNND5gierEe0RVn8cw7Rdr5IlaQEgU1fynvOf7C1
eh+tLxVqGs/L6Uy9n5Fk3kZDfNgHddwEep8BknhuDcFLSnq2ZOswqNtN69BZ409T5Ohn1XDNjbN9
t4igb7nvTCfYPoH8kXMgLdeq61Hbbe8sEjOXYjNblaT0HH2GJb9kGmeo7suqdhLQ1ljayKJdM2gw
XvyPAbswb54cqQQstgDLzdbUEJpF96Ckqb0Ye2sKPg/1UxLVpCPAkl1WRCu/okHAUDRv8jvcTO2E
xDkVTA+d9GkzuFsi5mp4lKNWq9OYsw879fyucrwaNzBFH0uRLj+yuakhmVWBqBAz7vsJv4M/MjnR
7fAq9UBYwzhI1QbgCuj7KO+poqPQd2LlHzgp7H+yfNTSK647U6CQvXMxzaaNhxNZrz0CVv/TNWQa
VGgw/eyqujujmnM/riIlXAVumTdAoRPsNeQo9xMfmzpvn7G9nE3/m+ggnqKQYyb6Z1usSet0inFP
NIJVfB+P+/yVZ1Hz89VR1Z5HTxUfPy8PC0kXKLjloCaFhTDqh9h4wU2STD6FsWg1Fu65Bkgr3EkI
DgbIdCKO+Rne4Do/OZxUjgySCF5BzJRhbzNE45nNKOCTfk1j2fIfjASYZKOYtCHhx9PLP5XYjdid
h/snaTopETt3XfNePehKuDknWW0FPuaRiLNJcXgmAWfKdnUatTZS8ts0KXa4L3tcX/qyH/waCLVf
eckZd5iMWeGBW6imXAj0ATG8K5I5JoJSCdrfqTth+eqDhKo+SUydJZs6NNBWzzjYUS0fwNVdU6v1
3h8eiosC5/LzIdwGhqgIpD3XBERdO4i/SiGcoxxewghFQoGg5JPasGFy5ixK8JYtGhuNncjGdhwq
DpVSDGfiBzO1+AF57JOcE7DW0wVUk9ANACmgZ7mxNfU4ZpEFybUGDY8GJdZtB+wkM0L7wnAZx0If
P5TkTl4No73iAaIqrwXX8yxmfa8v0BRchj2TSlcCorz7azlUl3SKkDuZ5ytiB6fO0PKzdHvVyzyS
cn+FoZ/p2mXXH8Z1LqaaRPekceUysPgKl0MQVOjpkpiH+5iTI6aEywRRh0DHZzEZehC6ydyLodwO
yrAfh1kP9k5VYW3JDfuzktalBPjSCbLNzq8NIUT1yIQgaerOCKnNH9hpTD1UC7BEseyaDS3u9wS6
rrnHnEDPCfgwQrFReI4k08m2d1vB7VNSL4XmaR0qhbgrkgHsBraTKwiXRWiLDsv+rNP7pL34O5O5
cjG0putKU1qKTlfOjqeeLolmnSUTy7ejDjlJpU+aD2Hn4AWzBejNMwYwdWihYE28eTw9bn5TDJ2V
6ntLwZstxYn+hDLjBkHHmKatOTALPw76649F/qsfJlUZlzGI2F3dUS0bChiRlWlaNsgIBjlR8/19
sO/IVE6wowa7ojLptGARDxa0o1gXYiKeh9kULYT70hF5w7dR2tvdzpeT3UddCANQYIT8TEE5Oqcy
Sh0iZxufWeCllLmYVt1cf2D19ohDIzRbGhR0vnF5iN8bV88U2rJZIwAWFgVP+HpzTuOH168vBjF2
Udsn/EXJEii6h8r8LHPCQuHHb4OwHewsUssimBBjsw5cCGO1qsAAiOwZ0BdzGyfEIy6vK5Qks4/K
n8ewmsUa0k/I+SS9ZoBcBpAJS+2BnW9Dvg/17wghjwg0Sm+CsdxBCMAf8Rxb/7zwpslQ741NHkfo
AqvVM8pKUeLcM75rX3e/B+wIZag1pwQioM0Brg0YfxpW/djXR4GKi4bWaQb7ZF/NK/0EZYtUSINi
is+eVrZBs+wghYQPZBCyet16IWNxtLAfsv1h6FipErIRDCCfXeT/XD1Zv7kBd9TqxDfmNQp3EU35
QBDLpckCZLc3SnqnfG+YY/xw0piLz1nQj72TixEL7g6jEZE3iN624EMJ4PBQSCcU69w11Yga6Pvf
kg7WhgOVhQbYDzzEjL/ZB4TrLWRW3MQdfMdH93PmcEoMuu9y+7IB+UY1lDnFPbNyghtxLf3HfbaN
MkwVA2CK9hp4ZM/kzm7k/TIv9+XTeABStu+1cwgSBVchrKGHSTp3C/dsEzdshzIWBU4F1aJgGrRv
nRn5V0ttiSC6cJVPZW6T9RKgHF9VpFe9m8/n6cqvkFY4ok18+Is9rTZrNR2/lXIr7JIDWDDmMkXr
7iweRevkEsViPbylBtzbFocwTHk3VSwx7atNwkejTftzr8+WV7GrMbPyYvod/o6lAkPf8Ho/Svz6
8vgpVeuESRh9iMyfCXSLo5Mk4U10mAFXXMi8YVVxR4dGjA5fsRG1Hp4AppG5/KOvW7Na7sdmF5Vv
rxSXljxxjcTRoobEPfFOfObCQEAMYB2OsE0xYaC04AH46C00EAIdnM5N4wLuf7hfRVOd54g7rsth
CkgyUN+2NZ4Xs1X+5Yh9sQB88GYntAIv+qqe9m0OWX2V3jmySt+Xv2ztgsW8+NdBoo+sBatrz+DZ
d07z93LJqBH7JIxd/i1BgeEfE5aSix8ClbaACG5cbA4cDslhKAHC9eSV7LsQYdcMYRabCamEXqdQ
VOdVLEWgS7NCVL2GDxhVHFYdWAKnbZUBpsTVtzcMTJhxRcg2jne6gPt+DENlUZZlc+1eX6lP2Nrm
/0S8rpow3dlr1bvK5Nwhw20TaICKN0cO582xkEmlKEEcZljEcQmb/6JTh/CbtItkeE0H9AbLXQ2I
2MSFFjzYdE4MO+ERfRdJrzNb/znj8bFND88erR391D0RzbHn3BwAwbApZUmbIZEw+MfOBRNrbt+a
g9oPAA+H5uBVTwqXVm9PRp0zUnWZaa/P2bbLaXllXHQI6md+0fPEiQiCTXZ4aGBM+58p8bAOo8tf
3QYcT8iJRWR9m+tuAINenTQXYN5l9MpvGM2gi1jF3GoRAhHLnFsAwNfwYQjZXdWEqYADsvmLJDGE
XUwKj7eKGozCT9ah3k5NKpzo+9SMuUpSKNbH0r0OzPi46lqwlM+7gy3+QOTFgaZ5zy4cCssEPYw4
QF3hSomvMaEawSIIkTCW2RpEGaYh3wXXrGl7YHPbTShSrxpRuRmL38sLJhtDsz3kXF/NH7u5T5J9
KhMsFF0l71S9Rik7D1+8LhHxHZU51ITbux4SrW7dZQ47xJ6LZdZVQAMyuL/XhutHhOHtgqMapo7u
NVX5W2GkWlZ9NAIHipyO+wp67mgPKywL85qQkuVobjwK28AQsfL3AbqdaTk9I2Kok5RQtAkqYCv9
chW/A+sOQ1nEiWwEPhgrui+zR+DEaDJrZ3mMUjP2xnJCPjDt/cPK6WChY6LsvzBHAw5NES6pyu0Q
F/h5Qgxp/m8E5WprTeoC+3GpBU+ZUWrLbCxmw2g+rbQxjMRcrWiqoNZO93CbB/s4n98Lfth4NeN9
kUKKVyAU7r2V25Vz4AiPaHCpEe7jEPo+JqetlYZYs+nTqcYZNtTnjOkptlSR8s6Z0RDhm+iv6Aju
o9fPbfTCgQNXngeNZkvcoav/lPRwhpqHIiUodfzVwtdwcK7LYPRZc26j5D6LAVo2zWcQhy94m6ix
7LoCgX7YCo3GlCKlPxjwTvfKB+7BP4Gri1WJKXXXsEP28mAAuV1w8JmHyBgscjxi89SnM2nvojk2
Wv5Ss86iRwv2khfAWAEKHmKFJw4+l/d8niaQ3J4YmFYwOpv7Kwt9v2YwRhTsPZMPjV2zN/C/wM6L
zPGVUFrvLIFtN1maR3uv3syJgVt/ypGdEfAU/SPaXeD54lUwQGc965RXoukCKMPbREQfJP1m0Sfj
ur/YKElTThxb/ElYtZsxiTd+Z9AM3HfyajAmq0Ee7SCGzY0qLD/1Nmc5dAVQP2qj7fJQw1LOCevm
A+ndQ+K3Z/dQT0hrs7O7f40nl1Y21BsSG9aZTPAK7DK0D2yMwV/hkwqtjdtKTU2Z6/9PLdwMGhG1
bPQfZUKAO+XzyeoRet1J1RCG1kcQJ398OIfEqllmr98iTzM/zfPFvb6JR9XDVVnDLkrpsoW8q4s7
VB5XVyvIIzXfR+/Ci2VD814wnOgXT257pr0c0Z3wQVyO8ASeaq8j9+sauEMM6vUG8qrLvJh7k4QK
rRKvR8ZXUnCEac9BZbvCWlHURcEHSXzUN7d76vmxmfpBL7GKAH/apWipo0N8N/aJ/fcDYeW33PxF
W7qEya/pl+PchFPwc/mIUUSXf6HLINackBX/Fqia9/tu8PnsX9ErhHJU/y8lo43QC7vlV4UIb4Sy
0AQ7D6I+4KyqnsT9xI1fN1tLwKatgg54ACWofZYYGDz5xu5SlRF4FEP+GBDBiLmWWcJUMfBlc2kj
pX9fB848csUQZrmEx7SHBkjOMbXbHpDvN0udATfybFw3uMIWvoSYgrDnowY4e605guey7LPA2F3d
1vbEgDulli+CQge5M3yLUEzY4BpoljTNJrUUAYmkcJdt/HQffEHG0frHco0eFBPwDuqhR1XDOgQo
8rU9mGWAeI3fmjroJG2GZWMq4HIycosAeDBX7tZY17BLLa9mHue7udJOymGzaxbAfVVd4Sa1glj4
n7YGG6d6gp6iuJE5aoqqamOs0d5OJwKN3KEWBpZdAod2y0gYh3HUhom7BtLixxQrDnbEMEHg6V2K
1L4n98BHwuFggwqDv/8XDsX+JTQqo7EWtMGml6XgS0ZI3CyNS2itwp694z/272JJ/RYY6DKf8gRG
dTfszTbC2Qk2HOicsgBHzN0VAupV0JIPFSWGf0b6cRuto3I1RJhkRFDWal9AhcY/2tkYP6B2wgOZ
Q5uweG0XKq4nZlhZ9+O/vV06IX3xF9jNBjIbNzfnTVLWWFOpI9DmcAuotKDm4ppJqsj45nejzGSt
0EV/sm/hWAnjLdP8zpSjdR3h1nrtawJWo6e+0C+uoiurwlkiT6lVxX0nHfky+Ym+jNr1R0bJkNwx
uhC4iR3QqQE9zTUTH5y2wi8/LZpIXH2drLQqxd67uD0KteNbA2hsfLJhoZttzk7jvQcH1g9DXHJ8
zNIF4J2piyjOmE+6L/EYcXYhfZ9dWHSeNrD+RQekRirGOFpREx+BT+Vhpr9EQT1JGmppyMZXS1YW
bXx7GYQPsLDqMgTQteOemBvUVKr5eftQOGjrDhV3sYt3yD0dp3wAVftV9n9zDMY5A3Yib6/NL2mP
8hPsaSRz43DTBeEKbKbKXqr6/bXLpDygwpKMeZ0/Z9HTfOBzqpSSYXa4VcCjnSOvBjzRPiNKvGo9
kStmUTQ2Tp/YGE+K6LS0ohX6qI6Oq09sno5M6CnCAGd0cE9fIXePouGnTdxESkNZbIH0AfCIX72h
Lz99H0ePwySIa2v7W02v3IdQC1bsSSgjK05u8ZpWkgwgvuk8KIEcpz1vKiNozGzSWcR3lj77c/UW
49TIinfL+IpMJjguETyrYoJ3m/RgvrxCWJxOURK3deKiCB542ZC3kE0wGW8GeGIcdJClW1T55Qpq
EijV1LzZ8c4vx999bARZqtkEGVIp1YWDny5FcMREAoEEPoW0GLX+QgBR3uRebxZDMTc8KuqpKjSF
GN9CFlI6QBpLL7CGtdElSndj94eJKkB7B1XDK7fTcgSR3V1Vb5KGphNy4Usdtt8ESpwKJTraRf2q
ymjEjfCJ7Foxq8AJGsWpPWdY/nMsw+nrZwFyMuXRWpTAkyhIJQUL25EknupdRgugBGudy9zBVQ+4
qOsQEXd6WoIENIexZItmKdW8eYuCh0mJPLuhwaGwvgtD4rf2fjNtGkPZ/5B6KPO6irqES+5RMC3u
V69KcGctwR9beGCD3e/kbwD77FVNGwpLTaEHmFVFMJAGFdBU62L337SdA7pxcxmYiMWBXbdPML9/
sbYwnEIUedxTVV68yM2Yb4QGUhAoNIwAquwsC3GpbZe++OUA8hN5y5Ijb3geWZHcLLmtlhY3Bs4q
+8AyQVusVeBnASYmrANugAKEQaLPGoSDxJj6GJWIvNaWTfOFNfTScpi2t/UU1hig7Q8YgrY2buBx
MArC8ZdBY3Dour/zccw7sVof3w2etnFR/RGJdsQ+UyP4GQQHLcg38pKkEuDoAt4Jl0IwmTCA7ste
k/avap9JxZ5M0Xz9z9xQ9MpuKyJzkHedOxgqpaeDeG+Qkap953UqRtX6BFeA+6a7/HGMEU+t6rsi
n/m+ZMGJKrbvftEX779EedzWs/E5dRnC5VFWn8eyNPWl3Dk8mtNfLkdwY9OrNg6tKRCF35/33jcv
imbkNnHJ8Pf9x98W7vPH3SzXO2hGJrKqdE3KkKe9fhDqhx+4V5LJpgHPYZ0lHBtyxn2qHYUkzXKO
UOYnrRT/OosJIL1L2eQkk0bXeanPrpQZC7XjG6qv49mb3ng9Ddx09OzHJxGftdqoAhmSMOB8zk+W
UDhSzMDl132QDFnHo5/bNXeVUJoMxhKid/TDinZDM0miWPnupjUHwArF17M0Tpf7KmWt3qdf8kEN
mrKBI9g4WTb/RAArA4qBzHxOTLDZvambjciRi/7eQ4yspdp0xX9B15/r9r5lsVAMSL/kDdHPtie3
IbwFgnORwoyrbpkwTBMXg1bacWj/w3waigWmrjgnEjdy07b358aKHsixVOqLKxELHyvJ/bKzj0Nu
ywwpzj2OHJVRnE6fZRVInUH44PN8HIdy3ZxlNSZTO7/PB24bXFfBz2+TsNBCeVS4a4tUF9ZGqoP3
HYGGvOcTImH6454wcNzx6duecKZvL3jstN0OyPg9n9BFX3CcXp35U7eyRf7ZwZWja/7+isMUutLa
xJRCfF+7Ctnk5tNJn42I3xj6bcD9BNVOxBIzkkXxajZu4Ol4dFuYGf2r9TxPDnEeiXgJBThyAGsc
lX7C1Ik9c+4La10DuLg+KVE7SY6H4QAwVQV/yhmZoUwYo37F6e59GBsjmr0x3VsdgjvJxr0uIIkE
si5J9tdcYOeilaSediRjWQs2rYN+AvZ/y9MHEMPZS7EJsMxqyW1jb0UqJEOtWyg8TL2LWRB9IcgM
/wjrxm09hmrFIkNERRAHhQjJEt1plAAliED4W/HsAWO6m1qCSRrGki01Jy3UXdFqjZr6q3l2/S1T
wuHM9PRg60HdzAvPYQOIk/PkwvYhz4txFW/8MbugvI1duKQZTdRgHiGrI0ZtKTvIzF9h1bWrjwcI
Ges0uerDbrZJso2E/X9HdLnFpeUl3e5Va5M09/UjvQbW6izWm4Pb7n++1K1was8KpPFbuLInclPs
Z2JLgryCWdzrXoA5KbjHUPiaeS8013RJP5ilrhS87XN/lS8dfJWZK1ItY1Ak+c1de7m+DM5/gfHI
JBHHrOgDIydqrMUZxrd6bNTOoQxKdsFXeOuebQKLZe2dnp7uXEHQM7S3LricTTJffJDS0n0IUJfb
1JaEEW0GJC06su5H45GhGKcu5d4Z+Vx3GHhBbTJmjtYAUhcste/Zebj+YFQ3oEc2SKVBYn06V+cA
tqcmhGGAJOzAYcIEhl+klSKz2+XGzvjEC8jwajhUgFHRLcP213Wnfd8gwMIE6hgxpD5UCgXTAsex
FEdjT7jwn2hH4fl1FpI2lySw1/MrRXohInSynWYU6ntxqXYoYMKbq8ksOHN6TgJ3TXKsGQ4fVVEG
p1QqY3Fcfk3San6IgBczoHlY+LQ2ctdZkqqmPLf2J4gzNrxONlK2VWcFsS5tz/w3Xujvx5zO8e3r
l8EUMxis7TKqw3lRuTFMRw0DRaV1RaTqFzmbQuG3RtQYC20TIl7P7YnVyYh3MnwyV2tl0iNQVY72
13hO11CWGbK7Efw1ndNQvSk1ytUJjaXw3regejcrA/KFmR3U1lSl7sZ/syVbwKupqhsJJpZ/Wb8D
beBARQBwAhBeD+sYmo2jSlG6LfrwIibw2yd5JvqNNo4wwvqrEjOloQWZ1W9mALFg4AyHP7cS99VR
tAZBsH1QODbXITLnqqEWvfEcQHYJcyqlo9Oe6jo0aPyGBIvDKRmA42ozpHb/cDdYCcfSwtyrzt2S
NgysSr3A7I/3rY2WekMg+NMFq1A2uZ67AkJfDnJa+sRj5ASE10POJkwWCTAVR8iCHzSY7YiE4rCW
m/syzSgvollJ4vQr88J/y3qUEy7E9Z4hSkAUxjPaqL0H8kXntLLpS0Y+HEVOkCKbmrkLDSgTYao+
cI02zyIesMffSJ39rGeecpuRzleGwztFZ9Ow1aYutRMOngXQHKTdIDF8CUE4om/NyJzcmtYMuJZ8
wJfSMHc1pnMEcRo0eqHUFCNTi+Qh3PLAdTTSXglbgvbpacpE9QcPFUD3R5uVCVfeP1Ri1te5r9gO
bE9ukLRYLgCsQSbR/RacZXo9QHAewq5cgO9B6Nwxso4TNAluPzRDyk/I/bQtPJKIu3zk5OwdlQkv
6Rzw6p5ty++nQDkAC+mXvNKolGtVNSxM/xVYCDZvw24kxUOflh0/WGPZBuz4wyN04v/Yg1vCRlyV
oQGBbgSAgaMSxpHhOMxDuUyV3xP3+V9ZWaVTnmGVVRqM2nSJIVzD3aSQIIo0FNKPLw0b0hXFApoD
xejVaH7Zw/FDTal/haHQMjHn+xyijJoXX1jBfcuV/c5LJ3K7CL4lt8D8Ws5tD9Je7lA2ZloCXECx
7W7XXATfDZsElxplTzht4pRD4Br1Eox6Agmm4AT9arVS7c013PHGNCbH4fMdGsyLaq1JuxXCSsSz
RfOwmbSIcX/ffv4p9NX33MfU9CuBmW0uYVaW1o00ZgfpplMaLEUvSYtLuT67+BHrbjXu0XnI7Pwb
d8pzxQOSMGi0O5hg48Dtpvbo47RFDwl0R2flKbZg/7elNDrqCETEOXxotgs1QMMKD2pbLJkbZ2RO
EP2dTdWVnLen3m4O/4gyDK5iwE0ZWdvt0EVKBvko//VXM93AoKK92eWbhDQJ/N+PMr2c/RYHxPBW
4SXPvazik2wTvKAwC/KuIzKXGGana2Bsbg7zZ41kg8q0TEU5AL8jMJBoSMy2b8udqEAyykfgxDqx
zzcILxfETNWSo7oDbxNCZezaCgjz8qit4SITUi14F8f3iXZ6k9LDtjA+OBT2U+mbbljZvg9fn/WR
yEP7reY2XpkwdwfRwoLHdMiqSZHYHcArqHlH3dqbgHPRFJpQooDgi1Iw4gEp79TW60p8TvlOa1Df
qzh7+vOfBbup0H3SKMnN9Toni3jw8IZDPHxUN4rR4xIr0PJzxw23s64xDnTCbrYFTRzqZHoTn88P
lgzfKmFC6GWeR2JAsTsrcq0kTkxLQAQBH6w7+T/EZf41s00po0rCr1zHdHPrHT8mHiJPC3z+Sirk
di8VuQGFbdc2FV1FA4Bzolt8qgUCgfwZq9Vud3Bu+eJoVEfrcwHoEV6z2QgLdfzRmzZx0yKG/1Dh
ZG0ezIo2JShP16WXiIMeZgQ7+7Wj46DSnI8kRy36n2ChwwVxt1koQEd/vGvLY4FgCdPHPqmpbG8J
zC0s0jAB67wsFCyd321kf6JEDbhhgXdwKZcUi6+CmOrQjy0QI4lyQ6cEfUWSC3XFdQo7y5SIVZ0Q
Z0bdyC5aWqANTRcvoSoJ1LDGMXN/qq2Dk/U7+jx1ySNvKea3BXogFeIi5EgMapjXmWYYND5MQ8FD
D49xuJYxNxLsrFHlq2AcZdv9EDODmOgZuCWDEXJE0t/qfjgovACvz+5C/mSvzKyCljLhtP0y0IZ7
0TBBP+7cKi1e62Fu7W8G4ATZwhwayoN8/VrjMgESn2vFTtmumPyxA3zHZYAt0S4V5ckGI/pNboey
7wBMPXibDDDCp9tKDFRzaBKAvmVJKqyriR+HYXPk9Z8apze6AYi15+H4QA187orFfD3rc5S2gcCS
xw7KSwhLGwpJbG+Izg/DjMAsYyDtHGLn25ki9Mwb+D6x2dwYoKcv0DyqhCKrgYvnohEeOTsAaJxg
GieA6gQxZ4rb5jbGtBa1C5WrAmmjQ/sRFRa6Lj4TD5yptTGb7YO2MECMuIVzjTAssmNtd+PrUgrd
ignZJu717wVTPaadsw51jg0zXY4lzaR+pJYDTYfqVKwevH+Efau88NtTZU8MPc3ZLRzlEj1Rwx0b
ba+B2B+egvVgZR2H+2hlJ6KzPP8vwvTeoAbzTSO1MuIpgbFetLRTuDnWk7/JwcfqQgS9j06ehTT+
BYGUo1gQaVhSqKhp0tZQdFinKXEs/+g9hKTjSlPNq7Ab7WdQLB9xkz5ClNhtOjiuUCLGpUTqZPnp
Rs9SHy2v0wwLP/DBJdHHi+dS1IbT1GmUueTUZmtFHUMyhgfINAj1L7udgbjOdni1XQwbQSWu/AaX
jBuFSH0xvyH33V3qHK3QR8nn1qUYr/J6ZXO9v26agUPmU2nJeyQTNa+IobNw/RUsGTeDHorzagoe
dcmAK7lRk/K/Kze/YZm7V21kotKPhQkWs0WHi0ByTA9MOCeUnh8Sl/jzosFdanQCibc7pj6fh48W
EprBv6NYnQIYIMUHLmd9YDz90c8WenmNy4SupxnloHM7Vw9WHOs/mvCRFjkR5b1JOIWK1yzvE8ak
g8bcT+/GqdAFw78/f7YXQZcgZ/vzZ9yv+rWEwtSctbQgbT95nuNKR8iODqwG/f1Bu+rXlNTreLbt
9URGmdoiIN9eJLxuCbpBKXUPvUhdiodgeiGYB12TWRbMHRuCvROvmvhsmQb5BQfzvFNJ0hF4d5Ld
EYvqamIoUFMhKxlS9l3VAJMXYhwR8jrhWp4LRgFNAXK2VEqQfOKAOAJVB5aKzTLhr2hajvC0ZID0
SZxocc4PTj0nAymdZeDAqd2SojX6ydYVbi9G/F8l0vfCeZxQMnZjo1I57HNIpWiiMr5Gw9kg5mnT
DGlnlKNxlkvoM/LErn/TFeP8qizGm0wu1NXzk63MCN6c6pNgW//OhSUGQCfJja9vPMkNQrDsvvlJ
Rto0nTPBzQ1FvxvWmmYIEbHrCUySINYfR+nuxy/izFM0emQOj56eSDD3tiSRxLqXRYDYoWakPP48
ZB+FErkmOqZ4tN2PmKkE6QxnqrXWLxrUi5BBpZFlckvtQv23ic7OdeKCH2obhsQebSYlTzw91qmY
M9Md2pSLJzRmbvyT9+4QgF1INEd+FgQ5XV/DurLGY9Nbp1RBQIn3Mzm0fhVVva6maj/Pe415dCwA
uBLdYzr5accmmksDQR6WO794g4prfL0Qa/kQ5UvthymOloUUE+HFGO+O3zRC4/1BKdwDKwnvVVzc
ds9teQ8fezEDgaYJa1jccIjZxwEZiHUr6xwBgjyIVTNyJ75GKV7OMtdGUEHLvWMfTvdoTnRN5jCA
rLWUELWm2+PHbnm04roAW05wjM7lXIvXa/9LdLUaC9S6xrIjK0pHmjjbHiJwv37FhD1k3oub36r9
eZZyg4z4Ci7AiOW7F3DgGoB1KKf4YK/wVPkjDJe58KFlTvS9SAOFbRvXSAwyMSZ1zMWwJFD2juig
60GBmGrhKmDkw+x6n+0fw2GbvDCWsyq62q8zIhaZNvmlFWsm1CyVvO8EI7T92QrKGtWS2kz+WhM6
Ln10YJgfD64Lf+Rgan7T3vveLTRbQY0bIUp7C6gtuNZXeXrPbAyMlmpPOdq7+5278M8gEZjOPD/G
cR2X/5njci9KtXcvKe/2qatokyvEh5Va1Yf3fmOMztPy7wxjuFAOgR66xBdyry9jjMhSjuspJN6L
btJQZU2T7uD6HnfbjepKyEkwrI4VmPbUtQ+5uzj7+ASdDLU85chQjQS6J9RG5xrVvRkHdtSzu2UU
WEBw+Cvn2/7b3B9Hk9476cVOU1Dz8f7CJdYdeMfmhRTWNSyH206a03A9aCv0+y93SowPQ4f2j/IU
0FCiN5LIQdsOs/Cy5DpJu2Gd9dhOkeu7+Y3Y/Yeby6Cs+A4tXZU3DSZNbWQqDH2LLDmbMOpPKXLb
Mdi8tenttsSIRnaRdpp/Msg3jpakhd31tAUpCeyPeQjxQcEh3G9VROrmaiT22d47j/giGpkMXgGa
DvUdt+rplz4WedSVP/Cski73OqgPZ/H7l6lcslktMNci7c4QcR6uYi/VI9E6+OPwUg25myCVHS7M
9Dte4J03N34qQLvMF67YjQnQwqVsardJitqs7ddTBUa/Lqga96rpuiSfVdbwWtOkw5zi6iQkVQh7
C8TFvilHhuF9WYgsB2r9lEZ09dxnhXoX5xl3waxlaoQPsQ7hjrnhSAkNTy6NwNvYts0NuKZ+bPQb
h/Q404KRxziGFEHeCtK8N4Ia1ESZwKDNhnUKgQQ7GgIb2GBc6KoLTvH903QaMRVkX6KhEPB1b9dm
Ieu/a/v30pyIxUXLZpF5lVu4xKTnmMC3ZXXetnTEIibscshFbZbYwPzwu994FhDhhrItxUjasl8v
3zev1fwQLKjB/BvvZEaibb48oNteXBO4dByWs/qVyzU7N2iatGxel14haaNU2dm2sb4zqKat39un
zsSf0VqSF8k6lH1wXf/N/mEtgaVHo0Aczj9HeuK4coxNr8zHqyt759+ovy/iylwAq8bX5HRFKWsB
4eTUW8xMo+SI2CHWgZ+LL6XNVMelfhgGdeRn2GiZidHsFkDlf3491iDCA0oCrzcQTrM01riW6s9W
kDwKkUidmOwO0HeyMnnIGpOyFF076/d4sMrrxFr2QsXqVBcXZoZVL+f2tcIbbRof3KD9xDLRt0oF
DhDgpKLeW40iRCYJ2AG/ihI02mayYyBn/sv8lJbOjlmzOYzqUieCq7Sc6qZ7RsqmNfPTeewrHbjU
uOFfAZWXjgmOyGeVkRh43BofKIQHRxjuUidmHbsLcPrueFl+tyUUKVrBVEPsHq9y6F2XTr5mr3Cv
x2pfDHwR3Lloq8TBeL6GBOB/Rtz8MOFDtoXNsnqkwDpE0YG1HMK9eS45tlt9VKYMN73SXwni7M5F
KAWTNcnyXnpjOZ5Vx3+EXxU4Rxih/Eu0xn3fMlDlZ54d2ZyNkJNtfk6KNMhB+RHclsgZy0A5N549
M7RO5GEjrKjSTB4t3j9UKhActF+5NKZ8iy3FLbWTESufBlUhM0+sA3+8IL5WlieTwsJIAoRWzP/1
eQamUBRjWwVNsN2+SzvzSXhpSwe8kRlcwoX+y7hquOoY2ULF7lNK1CBxkztoYgp2GPrLh7GUN4tv
lgTFQ7pRvAoowHb1U+enCzbayiJKx6ljgmVtVXErYsgPAu1TcieMohpFTKfv3gmCM3V24fT93wW9
+r2XFRVgMCSBWd4yyrjCZsaj3j+9+Lweg4rHTG00tTmAOq+72sIb0yAC3TuWZeRjfKJ2Xdqv9ap6
qmAF6acQ/OtRiVp0LrvKiVjp4APJhKrk5rxEdKdx7wfnZKgVn4I6H2mQcGxsL9rI9ZAf9lTaGlUq
a1/ZKifeoOBF8yGE62thFZbyi9lh7EeFin918HAjWlnno2hk3qDW2xYsATmk8n3z4GdTYk9mWbG/
wjXMeq1dNagFvfOQNt9BflD6CGepWFfnSnEAKpz0VDmCtDxYBf83wJpkhKrfnZcNEIgI5RN91HnY
TzmVX3Da8uvSHinO0MAA7w/uTCYBFuTFZ/xyOJSkUoURqPSAe4NNbHU0fD7uj0/HxXbaesGIHzzA
h/oCWFWN9f4mzjQuyaZUJGNkUkr3zgP+IkyKCdznwUG+MoBdgwdrkpuKPmczyHXUH7A2bAvm4bkC
+m+vTJUjRDU0Ojqm9FDSwBgIAI/rOGt9VSx8nOlnDJOrX0f7BgOWfwSY2bFf24+D+83cpOBZc+P2
1LXCHeouHO8XQW4f2Zt6ppujntwXqe2X5lxZhOdpuad36gVD7UFao0y6S6IJUI1+SyOyqydiuXxk
9GO4vlhpn0q5Z9t2Y0bm7XVjebpkEQxtfkRfmI72nXB3/+glGwvROnjKlr1cY1GpJZdZjyzXoO/X
z7ze0VzY/1mC0X32FXkKWPKXKh/N0Wvvc/M7PSUbhquu7104WPOdFpXQXAM9UZwDcYDId70qmYam
rp/j1OYhyIrwM25yzH5RNb8C6cE9TjatDc1xNY9cwAzJdaH+r3QpjJ7oCqX5T0BUbhLQ4E456a3N
mV1alrH99rpDXmQsi2lmorcCV3nrsg2Bmkts5DbCtikNxnaBtZPMbgPWVXTcvIrLr6M5jC6fJu7P
B4sDKnZnLbjthXD1Tt7ZvZ6zTu9nGvlCzrW4UYTFMRHN4SQv63Z6QeAZqTMVT5qGQ+qvYGQdtB2h
6g9VmV/6LchwV+mlBLPITlrqPmW8XBzjiVXWT7DvKgVjtLw9LP9925hhXI6gbaHCBvuQezPbfJnD
VZUjBWzwOZB/VXs/+/vC7OXuVYQ/Pq/Y+Ig+Ac5tUFlMzJcHrG7EeJwjQhIAwYG/533jF5WfWeDd
Kls3avgtJk32xu5Ub8YOMhr3C/Q9xeLcSLRpmxka9ZLyDgZcTX5ntW0w2zLZDdDA3rDQVm5Z75Yx
e12EiIA6hjMPiWhlPQF86GXIRT14HhYbo9Pub9A0BOeBxG1vtP+vTMEHfpcN9Jv7d3le4d0EgafL
c39bZyq6sFjRMG+SXVY5IAmwb5q3uURZwd7hkYptI3w4GVJCnyCu5hWd1UYOuXCb0q2SzF0WI26f
v0v/CKNpM6X89iCfR9uX1KLHWFUd8+QDTQ786mAZtnbiJRIae2fYaZ0pGAr27omdy4+pmmekSI0r
dIwMpxveFKOUfcBG/xxptEkieOJnbsXPtQ2zeEh9qEcYHFShNX12jBlxv2H26IakJqb92EgRN1Qp
ZxVpaaL4Z0WRK/idwdFiG3ZdF/xu2yu5gAQeH3F4UyFhJGAuxE49Lw5ARPD/IPk/tlrIWsdV0aFI
ts+0vrOOlTYyR+S30yLauOrCj0OeyDSfCJFmJJAkoPgaST343rUQL0tKYkRV6QVIgPIOllHq/Q8B
mBdOoHSuXw1q/FQtLS3pZknNt7eE+AbZTInmEtd5v793RbTmJXNiHnqSwtT1EepkVaa8HAS0Z7TV
Azg6sH42N/v8asaJdCG3QxBVLTZIdH6vwe13rKhOq91BHg6VFJBHs4Hs0Ufh1A/I26NicDctabUK
zAnz+SWUocmUggrgPGs6zCMX5m8SJ9OmlKA8qzInBkcFzBd4s+MsQvm8tkwtBqOeJUnWg2JStlpn
kdGjpfmPERNnwERJYh/ho3BFZdm5vy6KL1alHgmMk4hiIMhth9eh5NX4R/661xEK+4v9+bAiNKib
ZVquJlClmL49RIEfGlcQiY2uY9KWvvsxS7Lz2+3ZetRuFtF8jWKL0HsxU+Bc2E1E2sSQkcCofd5A
14/5u7BfqJ2L2SEIyFPnsISyYDvLhYjlQxJ6IO5E6QGDhHkTY4dv8QP1AFO9IuT79fmpPXRhdFg8
aLGMA8E3yMH6HtJVEqgi+f42oanLrUbJpssSXcyIjGSKChshndTwWB+vMDrQ9NUGMx3pcFhdzOTQ
WYukT71Vf8UtTP6zMrM3500pFrt9BjHx7trT3WPWgPwxmebNV/PXj8X2+qUW1xVP+JaO0MCJRG1S
S/LwRfiemq96GVIlnijogK/Oxt3PChaCOSSRF9auX8IKK9FaMdflsjw9DMQCIRU6I4JIL3yYoHOU
FkVpXFn35Xi7R6xnCDzmBrKicjYi60uv/JVJPh0vszKw+we/szzUyKRFPZzVJ3gMAJs8z2s22GNn
s7kYPNVZ1OGGOoMwHdJVp1aBrPF28QMel5ZepxGnf1JxLoaa03RMkZI+qtywMW9x6X77Dj3+89p0
3hvk53UymanGuRl60cENumnb8oe1f8ROsMOjzlnuDoWNp394/kcg66BdTL0iwT/m77DMRGULI3D0
5K2G8ueWpvV2xVmQXwLUAQuJQQNDcP/2vSvxx8CIO/zss0c9ZveDDIoy/Am2bveUnZmqXyzJg588
nvQhppTCVsKIuxFS/FZ1rBU89/G9vQ/xtIP6aQczJiHqr9hWaZPcyCeregyx//gPqaSau4EwRXXK
8zZldLoxtHXIXwMZd5DgYamkAB6QA8eb3aiGOmpJu9hwv1Wut/IYsE2IlsBHP7Ifjvy3pX9HlQaD
INRcZ1pJNODwigeg0sf/f/EABbb3TPbj/fgTxVREo1VsiqbIkzqqDTkbu/T1t/xAGaXwS5IKtKz6
v2H4qhA00RT7LB1+mKwlDuSRo3qAILNEkSNXgJGDao7+aMk7VuTEGgCph3f5ppQ3SaswUJRDJSmT
cU9bb85P2I2MwDGoNdWxJApGcqHLPERdjegcmuStELThn9Ra4zwmzqFBkrPnAmySE5sO8VS7yVxh
U5zU3K+94CJBrsa4KrdD2SBHT3TQiccTj8ejaGbrKrggtt/n2qOENXZVWxieDgBuTYcz7iXx3ana
JBrk8/2pte9EKseItfoE1x/+VBHjj7eZK3W1oGEjx80pQtuM/7V+uj8eOFW51GNpoNPhx2kBpR3J
huuZmhly6Rfl2p1wTzzO11rSjB8iSIEuKmXMAKcK/p5rLIzoiLICZggg/7EuVXPtf1iBTgzNThEM
kIIwPXH/+CuryT6X4BzUG45wgJBLX6CscEzQmQuabX+PLKsz+aAawrnIqMn8arHbd05wCrZim/3x
EZKRcv+Y8gw6+2CKWtctyCZm9q9ESaDZ+IUuHAVZ21gmYPgggWtR8NAynBlPCzzQZ0z5GZXW6sZQ
oIHtCQKxSbqQp/q24wCkUMJe0wpjvrIyXX16yw5MqW7lDVO4eEj+lpo6j9IHZHhRboyKkwE+C+pZ
pgUik/Dwf6/qUNJw+FSDCJWkq59dsf3Y9RnT3CsoBEg4vB/W5Fi444OW9529k/e887g19VZijllB
HbiG5WF/oaD/v+ftanvACg4/38KNP+txWgekhtXkJmUV2MLNoe18Se0S7+X3ZXgBxi7F5sSxHFoy
EmMtNEdEeFA3BCIL9WNf+s0pFB5+gfTpV7mjGk6b12ZKeNFUE5YKEqqLzKYnmolZO6YA6OxxCQYc
q+occl9Z3zBrZL82ryDgTNtD7d3AYN5oUoelTwWHYShf37TuTbrb/V7B37ntFPDUJwIesF+QfjGv
89MymIQYtFUMIBj3GA1rBgLE8Sjgrtdh8Qo0cRYjBUDs+C3EuENQ5HrNhviZHD82O93GRKu4/ZiL
//fBx7k+6+AwFp7lpvmZnHB/0vL2+NKUjyrK2rLsMrZBP/S5yhEtQK4fTcxHI1kg0XINQAWXFuVC
VzGdRApuXnlb1CJAVSpJSPA5Y40wSC42iP41dBdxrYNlxJNEo8JyXIn9kfIwQ5AUQVYiw8gd3R+A
c+v4C0Ey+1xW9u5XZyo6J/pidhV5r1Kv7a3DTBYBw9jm9lwuU2kBLqQRCIwYpQ5v5bpcuZIY5HB9
W3sR7vAYQAedyU6dRPt+K88c4mN1BUC4XqHhUrdsk3PkpCdg4d7cJb7wTY3VUdFjYEYc8PLkLbw2
cMvnhel8oznY3O7+3i4iKLZOhDoLjFlk0BHzWehjjmDJqLRvf1gt54Ss2HooM7Uo0O61xnP8/FsW
DVQEqCE+vduOV911gnwgaTn+wDyif+RlPvCGkHyMKde56wSjGauL8d2s3DkF+tTqoy91E5RlciAR
S8JPmCk1UnKJQ+TBWNg2vojdCspYQnJ6futXlE9XmE88EJiLKrLSG2eXk+QzBnMq5ir8CQ/yhhbY
OLaiCM+aMh0FFHrUEIsR3iKlcN2kytRaJizkGGjGzHGVJPx4jfJbXQRICM0YLvuHGp/EeeL3XHTs
IFfjTpiXT5JmZb2YlNarBTHnBtDt17vrq1xapBTgSlb+VF8qMAuMq6oPsXbzkFFmvbj6BGgyYCP0
pH08oNdwYxNciu8cxnUdp5B6QKCht1ZrEzAET4rbhu6FM8xLZa1S3FSgVWKNhN7a0CxGWaPeU1rx
nf6LNclkrU4Ys/P0zcIwu4jQDRztK5AvYFzdtnabJ1Af0S6aafHM6bAJ9ikY1Sy7QrafzSKTY5rI
XpHogUMPbbJ30zL8PjxcYX/gjtbBbRB0CJUmaBfIYw26XvjLtV7mzn6o84QNCqFch/YreGDE5JZq
mDebmJ2kc4C972tQWgYNK0gGfmT6ggMIyrdMuGZpSXUzyMGX828bbbXnldzKOQ85hNLj5jOFXks7
53xCSkAXopWD2qWMCYhvtbaXQIeBGzgf6YYb9dkk0zwT5SQiHQ6mMMudEYQnrury/n5jo7pIT2ei
AI7Zl6ZLB7qizn1YSFRQXYjOL82vCs8yRjU1lEqEfx4zoMN9Gd367RPEfoP2itv22Edqq2FjD/CE
j+9qQOTixn08PJXBAb7A26ecz1HyeaOo/QBUxPUtNR3ztVaW2N5vpQkXbmvyuH/+DLygTMQgpZGr
1g76mH786QKW+94STB5hTWEbYU87wyUA5YyTmWl0vV7qi0Jx1P2MZGqMBfVS0EuNfy6PXeQskwFj
VpZiVQRZL4GYcEQYQ0D0hDXBD5VxmbEpCcCUzIz2DklA3MQpM1+oeVM0RgXmytC7SMUIXFjrCjZ1
qMaJLpwnUryn+AnSGfmc61QGezWdRG7Lkc1SxaofO/ZFpwDzjt007ztd4gJWEnjTEAASklst2iiB
yeunP29plRvpZ74pq1bnnV/Y3Odc3hmZJSvvfrrK7GOC2Ka7Tfz3KAciQWeEijSLhQgCnllJA6mC
tURKhsIQTtzh7zEWVdSrmUTj6Tb6GROwxM332wn5aiTlZRyZzlGXIizWnOlAh9sQQuO+SGXpQoQ7
bC+chkQxn4IMJsvL/il2PVC5aRw9YCnSCpLuKkhhCANOtfrwOdh+CSd13P6FiPjzPizLsn6Lvs7B
vL7X6wFcHVaGvjlUW6104w9ACoWIzkELFzvtCmYYhK9Dt1J2shJdau+45ZkBFWMluuaW5gQkstn5
RzKMaKhFImM7xOXompvmkTjzeKaZ1gmmvB2yDpeEtc43dbpCArKpXddC0rbfDSbzcv1/3HH4T7HE
53B3K2DUH085/r77NjGy9IiaZc2banAsDyhJoN4Q1LGJI4MWaHdiMNQ7EOluetgyqrbPxqhOJG85
njMGvWqe3rwPbV8qhlFZTzN3kbEGgQ+Eeo+QatGSeb5LrVXiJKjzCRI4Cu29if3zracXr0s1wgdc
dEl7yLsz/jdaRZG40DZIKu7mdbgARUxsjOJcFlhSsLD0+3GXYSeho4YLzsDy3d91sOfkrzuFf4O7
r9xgMjBVHG6fzv1/NOcXgw/CaJn4dz5smY3Hfk9CREuyEHJEGelmOlSnkpe1ZQPGiVV4pATlxIF9
0uqhT6ECgS1X8FZfKer+ro9i/LFc47wEyXzSJ5RMzSkf0mmDFNzFJ0/dnyvAJzL/oYvhU2DTCxk8
5/I4/7keH2caXxddRjRH702QN50EtXL5MU6pnURvh8E/X+2kXUAoWaki3v/hKy0mX/Jd0kJAUaFO
YO+/3/EYv6mXXkKw9W0pn8SeQUN3iKDU72gXDt7otqAACZfK1gb77adxrJ2DUwfK83CKgQBhbpgr
Vj0q/c6lR/vwnYKGyoN/0OSJCQ99eLZAG9TGOf7YyOSiycS1D3AfW1gtnTwk/2DtaAJTMpjpTz3D
aGmZY9ObQqX4e3dC3emqEfl85qywSNzPJf0CCFUTfDwRl3sxW6YiD9jZ+2q37TH8XJd2IRSI42GG
19xMi601AKdMoyUDsGVQId9Rokz/CsdlpN4he2hvPscDW1EV/XMBGXnRc8cLEmNXijEvu0sF/rDV
mLOF++o6DM32rRVEmd5WNMimkL6XtoFHtG7D+lMeI7tsTvpD1KCEyXFuNHUL8nylwOQb5JT3DtWu
JJiIQu7eOFWFEYJsri3YnjKmYYncCsB73/PnEzP77tn0c+ZwX8DkYKALN8PBsI+FBhY4jUOmW950
o24eADaIGu4RJKFPqNiGURaXs6JEBCp0JQDY4KgnxPlX9aowCeBG6RKvjmEDAUAj7DkuHqqPCvR+
BcTnBq8AGJFeVsfX/W6VUqfKqEv+rvDasZNG7y4pD0WMx6+HKG722qBy2Lo6++ty2EtzTBWnZLWU
ZUNggqYIFHGIqkBDgSJAR9PWRFuXNvNBRaGijnCqYvuQLlWp1wJLreAHQMVta0g60wPeK1FCGtU1
O4pGqnYaJb30HyS4uGnED2Wbso5OCgLccTo5wSAIfj6dUP6Js2ObEFb5NIJ7AXmf1oywJnQdzAhH
Jfjqm0G8Mj8FWdQkLys9owjerVVBXOYKFB7yXWj5anuMWQOy/dc+MCiQwIOFgkduF2F2UaEK+rNR
Udfym9QF3zKzgBlEtiupEjTzH3DJO/AX/7uvEQij91tF5M5Nt2S62pU6X6im1d4Ex5s/6Bxxx7RM
oNYNgn6M0UWcLb4eSfEP5IXlA5xj8fdawmVdsUAdzn8VzkT4rAH/VMku9/rRT507p+TTGp4lzr8q
zwlfvly1jrEm3WnrcuEibfuaiAE8ZGxtDhTt/A2d35s9CFqwbrQUB6OKzM08VyBFd+r5HKF+LMKU
rkrdaSsjuF4b8xx8xXqKcP3TxRM690lgpXpzIE9lTUF8EaQTauLGWYKItXAWy90ZsiO6nrTtcbJB
7EIMFl3DbvSC9w0cZcyaKS+lZtydD8LvF6pJIIlTb29t17/KFGGqYiBzsPRsK7edmF/Mdy/YYe5V
quq1Vc7HUUyHlQoPwXgAG53UDb970AASRLQ48Bjtq7RMsc8mIKV+fDcSNMC0NRgQMHWOQMiJmBqn
JANhYJs/eKK3caR/XAp8QAmjrPOyAI+uPuDvZ/XOQVUVrLW6oi8HETVyCa03aRcx3CXNO9dP0OmM
9uNhypZe2BLjU4CLymmDOFbmNgr+8geLRQzgOuiDLXj930s6qMMMXENu1YkSvzVp89TUK26At+H/
ta2uNhhIOQKzCSmEvgLenlYLeuPPnDzZ8CVg1UEFqufsUiT2dlPik24D0dU7SRJCCO6HTu2Z+tfC
70jSVuHmYhl/z+slRcKdr0xo8WkwuqocczGgTA53IMekC4Lb8Mk9cDdWdTXRVo9lEY0RvDEF7DLG
Fq22mDB34lz2TcrPIv5uD5TTWRGZVPsyI4a2seDkqjnqVLLKIg+myS2Z0TSRuCNejjaYJZZ1Jmsg
WmKb+Vezd2Fs3We0YK8H72AL8/hNSuAdkMYETkxcWJlAzSxRBJD31AyqYBhotU6FXiDsvCX0Fpj9
WxBlGYQfhwR4FwdTGn5Fz90Zcq+hhiffLzGHF5+Bh2lHDKfclgfh161+WF3wBHJn9iyVuvTeA0Pi
90OeSrXopW/0PXNvYn1FDj28jA6wgqa3dVC9jfGhbQZyGDzHpi/QPm67UKeZpjAXBFnnvMouP+QW
dje5c1U9FWzPSbQ4AgfJlXLDkAL0QEqpUtZjzJloOqK7NM7jDqlYo3Iv2XajDm9AVi2Wg4KbFvM8
RUlXJOSogrUJKHlM76TeuvxDN0RxUckBPaWVLFC78rDmE5MBppHZrZfkR5GhQAErq8IuQfBnB1mU
eZHsrVGTBpvydbBMUodB22wLU+GD1OiUxzhsZVp1Rrb1XvBsVhdKa2oOnNf5XucQzhqqEF0q4aiS
didq1/buu1b3bZkiif13d9t0cVSlG5ABVIVMH3TRFNCPziTgpbf5UEjmUSRC1ZiLJLnj2vou4zPA
2ZACm63bRx0qWhdcBYb1LW6BfP8p83SSR9t84w8DE0XApcVdT8s34k2ZJzI4wZga/BQ4do0RSF7Y
h6WTaePIMXAr1nfHrBbKQ3+W8NDzm70P843bGZhnYgLQNFrufdO7AT3bm928J0LC8YaVMKBBKJqR
64a2WMiTN/LQq5HUwE54fhbc+JBwGK86WdBTTX+GbiezX2O++laca2nKyRnG/t1pMbz1CaXWd7hi
gSto5X83DjOufOXFBqBbAQTDYme0J1RuHPZDxkVeuw5ZN/WXwrSFQl1E1xD95Soabf+QaM4Ebaut
mKH/OGroOB4cvcBCg+Zga11ugnaz1F5gTRzQ9ALjbOrqnPUUNdpBvhV3+m3hqhd92zCCTdaAwxM/
ch/XXwpEMbiF/d0y0ZJa8vFRbm9xzKl0enuc6t8rUhzlQKe8+UU8e0ipNpS9cCImjbUxpcCw/hti
PwncRpkp46W5qxQPlnNkc9DahJ8X+o23Rn/ku9gQNJrudc9OxBAJG5+4Yiq4BCobNe1mrnpQYc8I
4kYHU61ZSg8h6oqOOQpY1cgjy4uhtNvg5VLpu34DRrt9q8xRlu5dqD5mLl412v09dJYwPS2TLc3D
6S1528NoFaAH65H5CdirwoW6523fFHx2EWEm7A3/D/gZKXRBPhax0CAaGQpQ1HUTQs2VXkupu84y
2JRyEHcpmu837QTRmdaT4PpuSGD6PBGX4vF3KHF9Wf/5D3X8B9dg0hXBmxVoc5pEsC1eB+qG8Rwf
/VuuyR8tnxLdP6iiSOJLbhuo5n2mLATD5kmC/HaOkdqu+H+hUOZCinBk2F1jNFw8nvijuym8TNMW
f3Bh6qwdNEqcC4P/PN2iUciWSfEIimQ6kN2uMmvuxvHe1Ek+V4MAi8+47J8hqdFMhAp2gmzyzp4S
Yfv9axRH8nyPeRpf4bev7mPPKnnOOVuX7qq300Im2zFfzX9W7hzacwcrxLVOIvDVnaDBzgTPtWCJ
K3YEgeCRRyRUO9ltLfgHH9UZNJzLgj4KYmMiai2pVCqQtqK8aNP3gENUtYeZ7XI4wVCVDhfb8Ppp
wzViSoqWnls9K3Zvek9oSwN2t7g47hJl3uV+easRHZOPPi2/GTN04Od4+e7aBwfCu0/3ZlB3Nt8R
sKxGgeIpM0YO+I1Nkaasa7GBl75lNGteEOZ+md2M9xC1I5Agu7AvOgLaUamStDXADWwMEoNuPEWl
vq1QHxoROfiaDCaJ9qrudxBNdWyvdnKpnL+frp7ZlrRah1TUDlUxoh+Gl4VzDzB12JbhW6ASiihB
w3Gwe2a9kZgKccrWQqkolcwi4N30Y20vuBn+X0VXN5PZScbH1eNE9dd0cQXh1vFjtiwKjscWvdPo
lW2FiuYR3QeMAiEjBU69keb+EoZnPF0JHKJp7hmWiZDKpcMbEiPqx2okUDnQ2nM9wgRkcD76uZ8i
UCFI600fsBkvcyiB55q4D3+rGz4dcyBffrb67kYZzlwHzzoZ5eOwof+JZWk+ckLGAAxj6in4PVk1
bnGv1pC2j9BZnOhjF1hJ7xHN5DQ5kzGjTXBiWZdy3AAeoKGuuMkyIZo//kE26s5x1piJZSt63bFA
5iWQF27ZhwxmxXnsb42isnArB2UklxDcGQM25aBrCIkPGg1P6ZbCr+TYIK3iON0/1uToJDy6AElF
5sgGaptsSG72idqpKrckJNz6PqTmyDpp4M1ThiWJXrPegwqEPBxwrxj+XBYJUCg2JthcaoNTTG7k
fXaO7INu4HVhPdiATuul0+3Nvi1n3hVmI9TKf7agyjBXTe7ahKV5HhAnpV6+F9qrgme2U3bJ7vG6
9AKALFJEt0z24VUQwqAzcE5WIHZEKGUqmhaihAG34ssstQx4qPP+iEBpT56DCyRPq09ff2bcYZyB
Baetym98iHseAkr1tMTXp3zlZXxKR+m7Th16O9OjR/GOlfU61OorNBUXPkdXZ/Ult4yzvLJmLkoY
j5c2mrqgbl3kdpOVbSXj+OqehgXV7IPLe6vFoZNf3AzAh4FTxH0baycjuR95d9Y+8k7SmGEOmSvm
f33M2vVNC6+piNmCHPnEgjEQHqkH1AgsnF+DMHkM1kUWZMSyXpiFzq1vDHcyiAvgF+tDnGk6hCwI
Vz1AZUDPVT4BxnUXHrk7UiHvRMQymr8TU6cgIN3e3J7eii9Bw3aEReDjJxGvu4iFi4mvbAvxIXag
U2pYWdfvXLWRxBjpYsIyy8/l/XzLez1dn9vQlb/8eGkmf+noPaBrgtCPGHvRm+poIEJI6OhZ9sni
JnrV47gUMGOe0Ac9gW3qJ7U+Yo3I1u6xjJ2kwOaxsc/ZcpbP9Hf92hx2lIJBtcWvStGMdiM6bDuq
cdph1ABi9dtGC57+bHyGV+PSsaCVfeYtj62del5g7mkL4CQbY2OWT1h4GjJk1M3jCNJWkN7Fg7Pk
gy4oPZzfCvg9FGf0uMqiJhiYasjk5ZOtfY+zraOjZeL+J8Bex9WlqRSDDquaEWi6Du+6fbEvNNRY
4lAtrk6vxyx7ll0aTeUkS7Sp5RBp6BXVqZmkyHYe0qJeJHYsc7GXa9aYXrTmB+gbOhZC+3uCOHQx
Ya5cLSOAF0d/GF0N06ffDiLNhLMPdxSB1mq3nDQgxbS8t6Z0r1kKJ7VXmUkX7oR9we/arrCZpPiY
Rro9VVbVb8z6Vu3Q1NLR7rr8OME6QBinBkAgdSKuYYBKD1wuEuF77xjiuzO3CPDlHwTg7zCB5Bfo
juWQhSe4LV6y3Rdp5rtyQUPxjeuv4xPzDlPlV2s3wt/nPXzkUiLxDQ1uhgLvxxehZV06IuNbpVHF
RVZWX+TLjVEYwx/ZsdUbK62/dw5QsiM5Quhfu3QHvCzBZOf7MXfdL+xG4MsFNycpwlf/uo+RMGNk
Ot+vN3yN141U8ftWrJW8eta3yNEJ/YqJtwxlJzGg3rKGzjoVE2Q5twFYfehs40N8g5vEf1u7ooxa
wJsYtdaOvtIfDzWQ4EPnPadXnCdJM0ag8oa/iyNedY8UXIDzujwFQaVFQyHVViVaLNrPARW3h9wk
eX/QdzyO8XfjESoSDGk9pllTsd4KcyyI3nHr9kSIo3EU04m/BUvaETYRwMHZu6ojtlmp2Q6yryXx
2kse7o8vTXNDmj94p0Qn3efl9sUIqRchxjaojO7EZR453YzUDwBJAIgG97F9HGJ9DirkbE6IrQD5
a/nDHXyuR9WPeHJw2Qpyw/yK+A5aKBUNBphvl04JRO4ID8FWS9uKJAIDrex+Z6ooQoJHnL82zBeI
wY9yY7fGFPvybJxU7gKx82i1h33NqYXPmZGBCRQuH7Bg1ZtZxsF5DYt4bBVXsWu4AyJhxNE+80UL
oyYkJ4cK2tKGj5q2Cb7W91elbyj652lA6Rzogm1yHu+yz1jDpQF+yoIlSnqgCrsF5QtI+DByp9xn
iULFXgPsRv5PsxY8mzeB4FFrN8zeVSJ/VLHfkijoMLYFflSf1amFv3DICnIjxpCmVp/d2rva43BV
y74OMLt6Dlw9Tc3SY/201JTc8MIFmlZ6sUgw5iAx5H8CpEvuY/iQBXPUMg073PD9njeqQmcHEbM1
FLPeR7iJr4ju7pJo2mTtVLV8fz2cWOebqc+zjvtAVkFdCJ2weUhPJ5XgDDLwTu7Pm3HuaI8ZcM4O
H4Fcku/aRdTkQ1c353oEBpHGosA+2FtDaXHMKC60wgdQoGVeMz4zisvd37dh7Tbny/K5/0Yxg9Ur
UQellf8GZo9v6sxcwY8ux7rCBVXNnibkpO0ctwr2srjjNLGUviqoW69fNNj36GzJ+SJCMyae513a
dtoOa3qXBxPSKrvAv17Oe4S27zVTqcTCAgQEDoY40A83CRSv94osDp3GWBHr8c4V3bys2B4Ipqtn
YykIa5dcfAU1wqclzefgZgVY1EKgK7vIcB1J5vsVSLyfnksDYKRauvE5eC26GwKv66wyDfKTsaHZ
+vh4yx3JRxF834xdJsEj/s3Z+fntjvJ1NCZkSMlW54o21twtev9dGq1yeIdVVdLpNpSw6P5X+IxJ
2e2Jxb/zMRyQgpfeuwXd4WabCXC4GW/5a58icEe43izVpUOSehY6ice7VntbliPucvsn18VRC4R8
3hIzvPEGpgILN3/YhzVRCh5pgL9FXdsp3vm+0RdGecoXeOg63qSO1X/UqExn6tv3R8KBgumqT6rm
AWeWOgt2Z99Tadof9EHptDheKTkuKu2s6a0IiP8TA8u4CzAFC9mNmbj6BqOR9gdowVlzoru+MTPZ
Qwk2s/k86A84xjLbavlIL6zCQq1zlyKap3+qev+SAsKUVDEqrJWxDib+M6ALa5IMwEZv9LeLLZp3
ZfdRevS4gWupWM3YwXGiX7PZXq99skCdMexE21H5uCHT92gRyr7SjMOBXDQA+N81zCYwttKLwP/v
KgIlDOFVSboKwgC9eiyyaYVeth+0x66s/TWxIc+UGXZ0JbxzdmUh6TxMyDTdXIes1IjDAG+NSnIH
Qb5c6lWGuKaA+Gk130J2UIrurGsrg3a3aqXiyT3n7JCBxW8FadYKxLjkSwhafb/mCCQW+ElH1ScH
NlnZexuA8BwW64wtN/Pdu+FjPLvB4ms765WLE5ZYILjGjiy0zTFSXRJqfKLjiljmB1t85g5VuGH7
lc5aE33scu/LvEeEdTCgzi+/wL1lvwzcmOoPMOy/DeIsJI37HvsRUJJVV0a012kUnq8/7ptaOTOa
pvz95V6Zb0x0tZj9ihldMhudMal1hWsf3OYv5UBfmBSZLZSJm8+A2NSevUPKdrkPeWSDg7FNlxLH
6PxPVFR9Wrszf7SPSiWltt2GoF6Zev6BD16OdJumvDGOm9PBcT7auISDQvHf/tkeJQAhkHMduIKX
S6uLUsKKCF5ynRn812rR/kzLxmi2cs/1D5GhxAw73jaVC5frObUMk6BIqqXAzyPo3uf8E9KWPuhK
1SbQ9Q6+JUtenoYPGab3rlXr8rGv0zok0UoJcREOQupMke5fTEQesj++y4HRe54380GVTHaaNcCD
pWklhOWTpD6vzhSM7qzE+PJQgzKSPdZu2LuPdc8ulnrP4VpbdgQci1IFTlBRrEVtqSfa57L8NcJN
/te5uld/X4dBpyQdDtW2l/ZWdVHVsJ2oWXVwnrMj4nbCL8hndXMylW8fIdVlAqejjcIU0fjhYo7+
Pn5U1iSaXAtdMYjseZd2cF/jVmzRm67XsUcG6BUoo1ueql0x5hJD82HIFVkdyGjxKdsKzFW9fX/R
KJoXjJGBYjMGfzt23kY53SytYRe/7tXjP2FuIGUXXLdtRU49MChwKwiZDDdQrXw4AVMoU6JE6hLF
OxknvpCXjr8O0tCL/P+jcZjDnK3BG2b6PMPOqYNOw5Pv1EDYpb+KZF4tgSHrUsiXnp+J/dNso9/Z
L0FJ4FEolyH+4fUUOMzikCrKj4TwE4LLlku5be651lhyQKdHwUSb9qVAJ6pxRQBzxqKRAnRgcczQ
TK0i66Hcz/knwzTkktLBFbMxjYJyDUoHCV9k0nQgNGRTaDvB/P8US5l8TnVo9z20q14TX43vgwqt
rOBgP8Cn6z5XTec2Rn4OuvR44YVTgolrhtZgsMvtq92/o9/arxZUCbnteAinudB1clv5GC8oiDQa
sv54X3QW9fkljrj5lWNU8qbM2pFBnLaFG/fhB+gv1WMf/0tEo6tJ7jBKP0Ki10MekYw5UfH1NYmz
G95Dpv54Ec1dahkoFiV1VvtT752PP5DK1s4QZmCyyTVshBB63qjkK4q5lNNbYr2xdGUp1dNbnf8U
0naKp6XA7KPcsDC5jAhhO9BjaOQYk7vO4QJ2+GYfrV6GoNiwH/VApX4PzVUQuYDrX8WyE5GMwH6x
v6bYRcq4MajBHul5lY5tABwCjtW+uqauhXjFDzkKxpBJIwPLdOQQdyoEXLh6YI8Btv9lziShfoyE
WqeJFM65gQkIXQEUePa4kUid3iUFTn8YKsM7QO8RBRECvJM8/xWKXG5c0XkLGdTvSsH4NdRR7wMi
KCMfdgWKFf98C+sbPCnnnQS22Xz+vxTs4L5l65UoIT+/9zsy6LSye3SYlqDdBY/4KYXZcRpqQIak
OmCvLz3vNXLkV3X88mZOSVjdjaIWEACXqUYevfniwqcwI6xGwMzcq3R8vcZNVgbdxilDMwyQFqR3
xKuCaYPK8cQ3HRzOg46jqJmpEAT+4+UnEccFAPSDj1x5X0E/ARj8VosLAh+ezuYkE6b4pYlf5H/o
I+J7LN9ZpKcdkZwzHb742keCeIvQcPWBJW7Lm5HJgr8CjvwQ5A3QD2bqgZs+yV0CJv88H7LtxGjO
CP+RYUsjGehY7IOqVyyLjowal3s7jKhJVeBAKGCgRxY34+AhP2YwLmC/gQhYt1gJ0zY5MSCEI9TT
1hv3nPIrCRfl7wDw1erSI4u8ZiKTjWq6Dloam1MLiL35sS1xCCcPEASuHGnj8zeMyIgKdHPEnJab
wPBa5ylL+zN8VmJDqyDW35tIvsf40bgkLfx0dZaMGMANZEJCGZDEOsAROrwfCWRPrvrRkSFMcM9X
vzcyQpaPcKh7tAsqyU3COXrTSDQNXEZeSjY+cS3iht1j35fXUokD7H0tXHu77tuMiLPvMv2LD4VA
IzQwTTb9xaXin0eB596mD2yUwegqtjMDjjAZLrRBdQx7KCeDZ0doZQ0iEBILGFgMHkiiTFtEDx3y
STvyqeG9k6QnqoyqSA1UA6vl5IdZZYmiojdlEXmGTTnDTr+ODhD9mBATv9aJYGqDkZy9hFovR+TJ
Bsnz4CD1S1rblEvq/Pja8lRzB1pE54rN+I9OSddTzkoLdO6itCVDF8rg80Xmur32gtvoWpwLvzbx
b1EP/2zWKVCc6d+SmSVjX1q491+8JYV7gThDDV8OR8YNEFvfqUsLaVZjpoHfqSBxlD51bV8uoMoh
umVGPSrCb/SkO9aT9JFpSCBdJptn/a1dBhUFAWS5Jkpmoxl9WxRQ5hVMCEyhfS9yfXyS2hK1KtFV
b6aoIxQjyuCzO36OXg2WNScHShGXMHEVLFvHrh7JfsxLXkyW+Fq7UJUdQwd9qH/pn5BvEdi9GHCZ
2gqSy9LO96X+Ez6yf+Vw+vNfUMk5ZJFr+AbUZkbGNoFIgJwgPxW+PP7MtxiZKZZqBrDWF7y4GLNT
OXj1XWVrfS1+udTaArJLsmYKGNUUhk1U6Jg9G/PCO7Vxh5QuszWQ+tGYoOD0KczJD25nydD7SiRe
AjHnoXia/+XdjXcgKQIG7wo41Lx8AITItbtiWfgip1sCaejfe8ck6iDmEXL9cjwdeN8sITPUBdE0
lsWLvTslLCPxn+6hDQ0N+Bd6aqpPLKOqY4/x5D+RbpGxkwxrE3+Xdxs70xmQ91m3w46U1Zm91K+W
fzAK0VlQOTbTTTRMYY21qLPRa3CSCEpuZSTCvaaH74tsQoLXuDb6BT7uBItax++LqYXdcyb8EuQX
fjtEAcWTVkpwehauaNT7ZwHviJ9fCmg8rFQZpEzAY92xnuLzCUWTy6wE0Euek5qwPnhNwdH5U9Ic
yZMG0wubfJIfMOPo/8Xy0oanaCyp8UtsV7SLqI370S3Z0eGABgvQnrPWmzwOq3w/lv5GYi4hBC6N
SAPaLkA7pod870fI6WfK0dWlURazVrDQeIO4+WaseE1zA/w0dQID3Rt9M3FXtd3s/j4X1WLpubE4
gij1V60lQJeaV1GQMZWzJtWNcW2E0KkVWbKes1pd81I1hPTJdizcCUt4XyvSrbJC8sLgCUrPXhSs
yiTW6pttTzgvVxZBp5TSwfuSDPuHsDABi+8d+2GerMSYSHeR8wAv3Dw5xe27sdMPlhQSbho3IipX
Z7P01+jFqCiKVItSmusNz2uA5bB3tk4aHzJlem9oATxqg5lEY0yX4ecyhKI3Kwlr6r+9B/HDcHOr
ag0Ocz9gJiRfPIRtxnDiUUVg+jd2WDAti9tCL7I1zFBydfG4adub/DqqSeRLJRy1LZNBP4r0AhpT
g+KGN3KV7OF8hjMBy6yLiB9oAxpcRMd2BR8XKOjgv/AA5eWIFVotDOoYBN3Er/YCe1zbv2F3NCTf
wkT9oae91T04ova0K6etuix0dAwceCd/M6FfN6GtKpPmQO69k016Fc66rOHOME2gGSlJ6RIQtQOT
LTM3JXpv240//0RWU2/sycxq6wmwE+YzQ677SQddJW6RMn8prtOwHsvMXvQmR5MlpqN2+fAio6CD
viPyr69s3xrDBlL7AblW38m3UYRWfwkwshPCb7B4WJOddczLE8GglzPHb7q6YUBa+N/GVe2+43B0
yf30HbFbTVyCHhCNx+EZGZv9utfBzzea/Rp9K76pNFFDcN8MCiREa1QxXugZJa3vCuUJA67S0d2z
9BExpOadLq4kX08Hhsk3sxHaNiThq3zKJ07bkUy1FYtj2KTVBN3cKsYxlBlexExWqq6y1WPu20gX
Eap2yiKV0xLUiQMg6A6fo3UgwmmSHaUrab90uM2BtO5KWT78xnLltcxnRQtf6TWjC/ZFV7fKYX/g
TcVFlntQy085XouoKm8vQIvJDaTuY7v7wusY9qYdjkL3GpHos0aUqKHxXJ36ad/rBUuJkSaS3xEP
iNFs3PiN2WwQkyCmBhExMJFdM6agoR16QLOhm6p9WRTfgNNFzYe1B2YXa5Bjwvc0cu8XY1imn28E
v3gb0M6LmmVC8TIueI2h3irYtWk52NvIDlkuOAqllI8QN3Iq6wlxqKBWZCejap4A2QS2h1lLCnFU
bfzSrXhNF5G2xoRoyvoyjeSw58z86k3qxoDuzxIJ3RnjKlrrzxOK4LmRh5bOtKQxSuMkJVDQMQyI
tB9NyisZbXfE241tabclvjZ7g3d932bJQVvJNm/FquMNNau+KT4JT+4J3kCNQFOtMY3iSEvqGeKY
0F9bVJfmkwfjye7wp/TLqnAlwJ8EhelQGUNTacKKSiGTf97gH9JY/bLBb9z8zT0zJzedcseRs/qg
P5jlL1wBXadulQDCo6QtQH15otCnXYejL79Vx2wplgSrFNskYLyvY2s600snQJqi2O9zQiZGn8Wo
nnAVI1fK0OJLTe49Yb3DuCefez2irID/lYMTAquTA3lTLUCFQuoaQJERhXnql43eT5bH8jXbphPd
a0pcUaazkWxHSwtohka7LqGOo+E7hoGBzXkjWUb8ULdmgCO0IbvfE5txk/3QGPHXXYsIjge4g5br
Hbk5X291Zl/gK39epaZNdyl4htqpgl2JqKDsKo0gTzwJp9i5XV5vUG8gQHSF33JPEVi49nU0eEnU
VwMYdHhTibMyneIameh9H1tHgwVh/YIpy5SolakiNHeBTvqjgX4AkswdPZp4lAmHcXWhHurW1Rz/
jDL0KmYVqHblfxIpII7uLrMiEugX//QASEPv0rcH99ZJMFLWjyQi2pgZeI2QeYsPBe2LGCu1knp3
Q+NYzF6RjiAk+Mg9FSejck3hvAAb5QF75QDzY14bhw0uLbwjgnYDFyT2/YeafbR9243gykcqNsmg
IFQo3eNoc4Zd2QMsAKdcWAJq5LsbtVio1brembZZcY5nYpRma7mcgOqUdH0QANqThYROcqoevn7s
yvQJ3nX9IIJGY/TaTNIHw7AmT/mOKQXYWHbvb7nklAiecC2j4rFHh6EL7QflhXpq8YaPpFQogGP7
AJaigSBYcTjS5kIKwZ5KIL+nGIaYZxfcWMZd8oU83iOYsoHQlIQpdYCd5RSR9KAFIUpR8iIcCW7G
YmIjAF8g0xKaAM9/JuUjRz7WBpTh9RYISbNba28pDuroDDW1iMxIE2Q3vhmAeFnIcimYUVCtOnKe
pn7UwGaOf6xJLnWvoQunutsBb1ugBaKvEJlCji9oY51lukf6p+EjiUyiyWbuRJcIRpci6cNZ1bwS
NLBK1p+2uS1UEaWbDcneWhTTuX/sa1Ru11lC2YFoaD94boUc/79EECeWH0v9iyWEM7//dhc+/iIr
D0ueA2cK8spB3u7DlaHdYOLgYf0XqEk9sG/RfJHJFko1XrNUok8ZWi+oV+teFoVQ/yy4uCsIPXt+
x5ksP6ykpIA1/etN1lPm4A6YSlnlbxTgjleXxpAwQ5zJR/U0mNe82ufx/ZiFBiWGTce00oyZNlRe
kFLE6pbTbzO94oJcfTO9BSeCqCx3+F+3XOjp42FW3zNytYu2j9zJ6nrAYOagoiW5zmHdmRLsYdpY
ohgCkOGD2vbbaXmGjtysSD+3P5O9Rl3hsV6tuKYpa72zL3Nm81lbzDCfcW23IcpeRhrM5sWNNDo6
VV5qusTbEBEGj91++QByHyZeoNmrTvAhYRmAzkk7XRMKKMsaPWzF5HPvZx0NEeP/dEyosCfO3deA
BNOllUmANyN+6I2mr4DSvppsH+N38YtuROZmcF9oqamtaUtvwrI3lWp72Xm76bkhsROHil7ZwxnG
93R32xZBuVk68fh2x+p2PO6uysQZbp8HYGy9p8DpbcbdlDI7W0XEyLp0zepsm05RtgU/6xPkHbZb
PcLAcweGLdehNCP73zv6CkTfS8t903vBH5cXdEnQunxZEnE5JhET0oJxh++g4Q6mrjNtGNUmzddT
jtcew4rEuDD0e9N4NrDsy8sl7p2pPV0Qb/NVmDtItxkR8lHN6Zu1DSWje1W7wDwCXEXvgY5VxQCG
Nsof2Fov+ZhY4eXPtyDLZ/WX7426JkM1Ga7rRL9ipLsJgq5G97sqNy+ndzteS+BkA1vFk2ZaDZNj
JzrYC5Z1xx+jJjdec21EtqD9sj3ONGsN7nQVXSkgURAWcz9uPwA4Y3HVwjcURXRplGvM5eT23Awu
gglb4Z621A8D6ZQcE8DNZ/aM/Kpa2s0QSdux6JRCfbSt+In9AVvcSgywevNlgVqkXZJztmt8GXd1
wpEGkC3eSeQJbm9vEFQg0eFj20xXH1IM3H6DbI6uzr18KArRIa0pJQgmEDYiELOs0H/qODrp3rQp
xYAv45kyOX9h04OICBqokuj69Vqry1fSoAvmXANg3aMsw7EgarXHFOgT+2Smks/sDG1gCtK9uPJe
fbu2SMNNqakuJNc2iG9FL/wRO/7n5m/KeI72NeSsQ3jzhr1mHnYWQhn9Uez9U/UXAadzqNz1k4Xz
bbR/jCChmcIWu9Du6i3zeb8OqSwSHnk/KWjlTHbw+qnPQFQT8kjyXHCLN6+j6iF6YlIi9gECglRx
MTGlEqWoXjo2oLDXMmJmYdfWBJvTQbzk1aEZVUZKFNcrETfIIXSent+2QBNzExYcZg2N2/1yjlqK
hn1mcrSFEftDwh7qrHTOXYiKbSsSo2TXIsI4aYROg5hsqW/eZBLRgDSA6FYXTlsrZ1Qt8ZzRzkv2
qMBQHxEC0YDfGC3HiMZvqZGoePDR79Da18lqvnLsS1Rqg45SMUAzn9zaGZX0d0ojCWxk0FOX7K7K
h2q+/SbUIBRS+tp4/O1HC7YYCkK1vcauXlcXRNvkCo2TDALYo/gb//vTSLLwZ9dxkkvZlWp3zzy8
YCfHehEwxLaZyyl8DE/62N7JQzTO+7KxknNhj9Dd+2HeCDeC3K/dkwcaAz7K+qmtkihJbUpMnDOj
hsMT9pO/uoZJajcl0u4dmkqj6PvbU5oFyIe/PcHia03btP1UO44fvG9K0Ibzt5JYqwe2bh5KfiHw
D3vuZPBvdm87E5MAYHmpWppZKkh4zVhygLV4uJW9cCrkLZgsMTi8fySU+oxfaphwLyENCrhHgRVT
jE2HhlmySzZ0Sc4qoZw0TulbBIWBKkHHIc9fbzqQnH9Bgbut4iH/1m2q156YJ8XQt2T/5Fk24aQy
+G5z+6kio/NHC5HhKWT+8fz5mfxMhiGtj/0WiYczib/vWsZ00ieLeR488VPQpCjwUiqSAs3flSLK
HP8l/oi+ZBu3WKbmUgINJXYa+CKBBhIpOsNb3nZMgq4kyC/P11WohMrB5R0istGMozZvpQdNnJfO
wIk8hiYhlZ6jE0qNHj4LVhtab1jL0KipobDayee1MD/9xV7gQE7L9Tmkin7kipXy/RSsX5YS0Jgm
SjqcHw0u0UktkIy6+CuJ0ydqdOPvIdUVAIA66RBL4fhF625Tog2OVHWV5+H4FNVbFeJulPyIRg1v
Ow8cYl3y3oNGzYCbAtH8TsM6g+qzQtICMHEmet2q6DCWrQ4uq7wuClhoYUYiB9hdjIENsJzajc0s
E5ikm38Hfd5ONHpeJgTR3KRZy2rRqy99iSNCjvvKqqfL9nL88AmwYRUdbGWl5nc0aI5Gj4OhnZps
r84XZjg8LyG1i3KE6iGWhzu68EdHX+njawMndhS4YdyJDnmOfJSZ4Cu190g1ngn+24awU6++7xDu
XVw6C3JzcFVBXCeND6psgs2wwFqBMHKOxlNOI3ST7s/fwdKiWsp4cl5u/ZCfahEE9I3virR5BOKj
BSnWdqsUKpsTSj9MXqNg9V/b/epUjXnFy5XohuxtkuYWGDsi2IdMgiCMHZ8WqacO4DDcisJecsKX
df9ohh29jUeUcXT7MYrKae19Bb1im9DD3HCoLhppM3ev3MQjVyZ69vfpfjDXIkDzHtAnXhPGZsob
9p4EswXW83dSxDJ4Xma2YVsLk4dNn+QJFyGboIbeJ4oPjBlitjRNPktjHoXz4/c8cCe7Pq0JRzW4
TSvHAOaJZ8yroIu/CrdxP8U1buIk5vewFbQyzU1F/kbhZVFY0I8NYYiXQCCEG/H0HQKE3aFJ8/MC
N11+VB6UxxP9Z27elU1yp1ZA+aNkUxTM9ZoV440nbuod1raRJWwS9vWPVK5MPlFmmz6wNlnFKViR
A+rkpXQPfP38fcI3667ULmDRlyBBydnOAIVs9AvMEOfiJxq3Uf8C9JkBgghZD96LHpfTvyGgC+hI
vFETjyxKJAr4Ul1G1JGA2N/mzmgwDiU0W+uTebm8l5dXtqrNXgFN9i84aDpbsjBLJsmu6W0pgIA8
chmN1lrKGPIneviDZlsUFlxMQUTd8XRXsHFpkZVsTQpiMrQpCxMOnUoEVnC2SQPPJO29qsyqZBZd
FrQm1aow5UUgGFnasfUfxxMUueyVZSUWvFgG+dk1LNzoZ9fpFITz+p8XYKHJPODZPHR9LPIAeQIj
XM5egeKZOpSYbSRTe2nzC5IyR4RscPmZbZ7TWwPAEs1HXbMfu5uKQswB94hJZCJpqaGySodR1WwX
cFb5aFFas8G2Cr2pF7+MbNpIZ2WtKvdB5daY7mE/eWeYXAk6PuG38zEwc0qRjNaJGQLp9puIQhmC
jhGGSXGo1GdC03FTR/cNhEUwrshZpYqIBOgXRmo1MxnvVBYt2/iRD++mgBOcoUvvY8VjjITbk7Fn
RGKXZ5GF/TgCqWy7/QEp3G9knphK73ww/0ehP7dxBZCQGk0YBiyU0/cFXpWdM8oMOpepq8J+gKaU
Qyv57IhzIGLJY10GEZGI2JqJSW8rxRZjlrAs8uEdxEG7SRbS6egAPQ+hh5nE3BdFzZD1iO8XOIwi
51ltcJ+mBTV0yZQVmy5lODNEwq6Z6676hFn1AsaPog3qdpvN9r6bxi7JLfVq5G9rwF9plhPd+UOF
8c68FL2vOjNnQJUuYMSkTzfh2NCKHO+0RkbYCL3+xwuJ8K8zmAXdPi6RHPIYFd/8JQd3zwaUiP77
05vq3oVgAVvERFf34qIInxgwV0iOFwFoPMU8rm+P+j0HVIlZH8Fs39bH7LD+RZEs9yFwQTo80+Wt
5MyDfqv2vDh6R2dvR9vmXUaI62meOms/+PPQwFbmp8OlAcans0Ix7TRtMwbaUXAgb2L+kOGayoZ7
7vvL4mnibFcJFQa2jy74r6XfxIONPcQDinoBgaewp9V9yWj3J677QrIK7E4SOWtBeLc5DxeyYA9G
TnB8OuBLJIWri2KFYogyROiZLBxTlU8Jj882TqWFOmt2kcHd0w/2o0Bf1EELLFXgKuGDbKRvF/Aq
FEUeQ4khBWrEHyqUem06wuvYk8SCPNAysjiyONidgemELuS9640eFISiE1f3irpSFas8OtEUaFUC
NT9IFpNV5sbR/jAcZrJ4XuQmILpueK5DGkmilxXeFbSMLaS+6GkffCCxP+p1K9IXvd//jVlk2ONS
ZjzW+d4e0jXJeAJ4Rkg5DH1XO/HtJ7YLpes17vVhFGnRGd7uE3giW4VKBOFT8kRK9xOgOQrsNhcT
gHKFxZcpJ1D//M3V7E0ovjNcIRG/x/KIpdbNIBYfgFgoQnXFoyGZvcoWI5jyvIpKrE96Qcq6ItIo
edBcx7eKxr5P4cNQ04GxCl/9IYF91opDQ6aP2QUdSud0Q4kOPJDnLjzD0eaT+W+qVx3+Nj1QA7Fm
uPqBlEbz+UZcWGCOjq9G1i4qQHeAHi2HMpepvW/Q9eNbS4eq0Qb0IhZV0k7JX47n4PcNqk93fr3m
ZV3NJwW5F/nm2VD2Y2U/q0hXKU5Az1TXmI/b0Xq1kskvfzXO/cjgZi5ZqHb10Iylfp/X+o20CQcj
zJso0IdEMGCSsS0sT5X0Q23NkaC34FKk4dnhnk4GD8aVNwZ2kiV5q7SKbElCuPD8CNjzr/VDAvrw
+jgh85qmiX8q3C4bJVs9Dk+/Dc4Q14AqsHog92Amkin03rBT/ITITKjW2vGcOP7TvunkJ5MqHu8A
N1uLeXnKWjdmIDhqe4lZD/T3VbGejFTI5fcmjXdGFUDnSQlgAqn3J159C55XQTwQJruWzC9udovJ
NWVEfN90b/JCnM20cz+FQKBmzy5oJZVmekaUFzuqbqO9hDBE8x/AMz/4g/Eao7DwNnKVWRg3iyyA
DKLgVt86RlOvnbyKsrGi3jcmwn1/Nui3FCQt3H+yjwVuNoBsbB5hXgHZyoUd/J23MPLTjbvYI6WZ
TuUzETFyRL9Om1Cpm4v86Jbr0A60UF4L1cjkOgGaVxwFdsK0ZjwTG0JE9JjxlmRuG7T0XEKTtd12
lJjaoYsdcQbxv5lVCrdx4zGvl/8/pRxAyLX/unYwELTxCS1BothavQ5b+pN8f9+wXXdTxZgrNd6x
bs5zsNdEI3UKKrLzTfwqH77IpNTKCoGnBDMSbUKkEIqJKMyyfq/BnyBdw7M405t+ACHuJyPobW7+
YJ/d4WRQQi1O/1YELOZQytHQ3bwAy0YEb3WwF6vJ2yKfAuNbNDNbgT5058/avLEdP4lUdXjh0avM
vPAnrbVz1UzoSCtNFUtcK4XnNedObWzenLkXrIGzh1M3wZG4iWcQD8W5lRwdgcBMzIjTpROhKFYj
wsO0mH4I4C9018nr8vgv0hNXIBpm2m6tK7+9fCF0oHKJl5piSlj/mig2d36VVOxiwMMnxAcFvUew
skhQYZJMbXOfhkqiP3yV1g3tAg+u1/NzTU4FuvTTXN8kaFZC1a/WW151DeGdIXKVSt0uP1ts6Qpz
X8jEgCENFk8H/Ff6AyfTGERSMHjRQ1lMovSAWnCD2+M8I/uWzthExAb238QQrwwUxz13CJ1SnXPB
6mLc9tfsUKOzXqIkrsjF+z4Q3AU89gpU5tRm4SVXEqMmv6Cwt4mQpGo6cHo58uY7MjDWV2EftSni
LFLO0k9vj5869fhwO2x5VO5+rEzMv8G9LagMMTq48z6N24Iphs7bCNfV4C0aHWntHRdjAbuOu1oR
BwkbgwZLWD1dgsC7OHH9yditd6xMIrtPMTsSjcaE9Ak3FZ6cd0bUbLJQ9itzXWNYeZ/Jxk6w8UPf
QJkg8/xZgsa0PsNf/qfkW3OlZy1XiO1IkvZoQWC470s/EnPJhQRbQo88NKkyxuzWp3HMITzPGoKU
nyKryYjw/4trZZUhjR0HGxxZHpBZNKCCipWGMtXX/G3s0+VU/UWqtHFtwlz4tVGn51mSHj0Mjc24
4XIxVyW0LxevlPuJ+prcC88c9FITTRspDxUJsQZVMtJETb17l/YM9DsEI9xxTLAGWOQNjDxsxbCO
WcQ4fV43hItMEj5l2DMg4kzF+iGl4lnwpWc+6NRiVgRi8t4U7UOBZ99BBljX9nf4Lwl9BIzWETgP
CH5X39AnGx1ovEFeKMIVzZd/52NDKXIPj3fWJbCwTRhbddVuEUbuzYhl8Lk4Jhr2Aq9DDniLXAd8
3FkDcSaB4eaw5Ds+wm59cdSDGV653aiHxAO5o0n+4BXrhIBITdCIo61Mj5NiWsdFMt3iLHA2OkT/
J6rrBm9KMo162QDn+oxDW4scWpeDxyWdU1tXSfrDlL6Kkxj/CZALAhO3pfXzR9obbNFZ7mfPO4+k
IM8xHfrgR9j3rsP21ZSp9NGCxaPXJ0JDNWnho2pkBgmX9O58R2CgpJsWiQZ36UZUu41qKsIfdYgr
bw0aXyHDSXfY5FvkMheum1NBUefBQ8UTtd0j3aXkCI1mpWABebElqtuFZFq39TMsJ62NHrbRlC5u
oB3bvC+02rMVvMyuJ87bu+WDOPi1ChM/ewdSoNR3b2W4M9RFPDAVNqPNHikdVHRQvyMrBCL7vIHj
hGjQ5zvzA5WRpNKiiBSZ3hV08LCTJJl6GQp8In/Q7isnf4Q4KGCp8Nd4oIlHWR/TLnW03JmQsirT
MHADd2FvHBuAogFuc/QCQIbIzD9VHqLMkIXaw2VkkY3hAVc2pNz10vwGFwcC4wmNy6hBYNi0EXXW
WJx4naE51oUNBh6ln65m1O2pQlJl4Odzw5ws4hHJqRXkQ347jF6wbEyBz9KNcYXW/qRSBS2kmxHZ
OYzLQvPuRlnJyLTBDMJ6ioWbouJC4l1YiIeU3NURcj7tSpDH9eU522uENS1HpFUwDeCKvxpJ5U3x
YIppEMSIOFYu2hZqyxYO3THkSdS+o40ADrt3K4b0OfV7DDeuHBnYLj2MGnWNj1E6Er0UwGtatT/k
g/9N8cvnHfu9t+x1xzESagIgbyvFSmAY/g4l9GaiJ9FP0uEgcbzglQqqHSVnXnTLWzsZBMkp46X5
AuXLuLl7u6s7+YcZDdwVDMyEFzPW5nDZsf5liaT3vgBi4x2Euqfdam1sU+qj9p4e5Zu/0S8yXLNB
LEANIDYjgz+5BD9zR66sHcDav56KZJJcQGvOuMxOb8awWkVVtQPgxD9qnHTvHoK9u2QNHikU5oGS
6tFxoTm6QtFO/2lo9MbK3WRV0a71ognVmiHsGUb3Lb6BrdTnWR7yPB3Wjwh1LynVi6MU7p5bq1PA
EYrAiczqfjmTFV1IijJYogHWT3Ld15dO9V9TQJ4vy9no7f78aK14sOPO++wPywMQlKuGSo6PEtxx
1YKzis7lwJ/8VQbTgFDa4FjHiMoz2Fb6pkkSAaA0cxXe0u34XQmR06y0oTWiz/tZl3SWdi2Rb0tq
/TsLps3n8+ndQbCBLtG+rWlKxM/xr+eBkmGh1FjuwNSHyHtHai/xor9HpnjDr3CDX2yIxsIRtsu/
yy7hIoiusCxl/t9IPmNMLdgHWH4FCEjUYhkC33Ls/vm5SdXxLQwMDLT1tSQkS8UEvcsc3oa1hkyO
F4NfDDWMkHPvmf3cG9DgXxRwHXTKtlLEk++1VdtE5cb0j13FbGwl/2veqXB2MvONtuGKBeAwNg0I
kAIbHMAYD99Lao7VPGLjpgn3RM7el+mp/wq3QopCf9mTCOTHdJY3Si8UNb6bJ9tWtI33P+PyzVmS
5UeLdxeJ2b4nNC79/ZmbB3X+T8Qhp3hyPeYTko/AYRFEGnIIEdaCm3O3UjYq2xk/fULRlPveuJLy
7SdzVfqzgj1etP8RNw6OdBo0MXITLA2eaCYX+ffbGcnz2nPwMRwqRj4NtXSblDmKDWsBDrrAj37d
dzvaHHln2AXwbj8B4ZR7ucu4PKafyhRNXbZmBJygBhRmyOzXwP8w7dzRBL4x+jb+b8RSXtJ3Mx3L
M/n2UgWb1NrWFuoG2QA0Ze03cHxyn+JRQrnK3XvD0CgCiun1KYg6FHmgWjp37HYVG1y/VaBTxWDf
VWL8ERdjFVHvQDKGP3j4+AviuHlkFsvOFSbtlGxNoWnC2qmHp0AWTU5iAYtxlZWkKuywZ7xvOV7S
1a7ebwhMttATAQQ6SpnMmZiisjq3cTjQJLlpH8gtHt6/mu8mF1THV+3Rmp5WUfXw9+y2GHD8InGn
3KIanzKcVRhEQ/aT/E41+kKv1sc9cC/3vea5eyIkLHGud4QnxPKGoRHW+uClSIeomUhLELVkZFbZ
rQMmG8/IVJCfI+DwPHxbDm0qMB4BMf5s9s2AcUR9Gn0P4b/nWHSH6nyxhA8KzRFwk3bHHY4jHBTH
DzfEISW/TPQNsfoono1UjdUd2S0vm8M5W78ZLWWGHjP1STDOVdONMhy7mtw+M0Bn3xTEjN7W++HY
f/QtGRzVVFbvJz+Mgx4tYrevYXHlqa1hGvTlybORkamTClbUQyN20ni9CbGh8UF+0IKjOzHm9uad
vOhHY9j3w14l7ey9P2HYxvqK4VAMK05xmgYAyJ9DDIB2ZV1yQzyjwttA7K8nLj2n+tOiv3YAxpzB
s7SBvioROjnpj10hI0cRF7ut7uVe6NeABoA2FLQQezaOsxmPoYELGUFnHZPky+P+hFGBuHAtRkyL
dSEmQNDl6EE2G+F1Wp8LzzmlBhutD2HyhzI6ytP0zyEHhGqiu4kHHjaPbIor8V9Mk5hScnErBaqy
MrclcXi6O2wJfixVF8AieqH1/ymrjdDX1U7RqAe7Zm8AlS7T+qh3jF3KTnQxagq4RTR1AmGrVdJE
/aiGhE41WsmzeaFQGwndxU5v8EIPSAzWLqtb4ITNmTaHS71CqV2KWznQfQCkml6qorFBY85Hy8df
L6jk731PrCU75s32aXeDF9SeL2vDL3Ccj8c2OZJ8MNMvFmgEFgKP9Mv9S6RkBOSJXLBmmpWwtoOQ
sr5sMv1RdxFOs4yRxIY66xfTs060SZMWezWlMSbj8VdDLzpU1A7MEwUgPCHY/ZqEnqNCarDSW0bo
wLah6HUhk54csK8eyQD+2pyoV9BqVk17yfx59WNsB9TWXnAPl/M5DEQ46WHxlWDLBT4JUCD3BsUL
P2g3VDa1cY0uZGKEzBVOo7ClP0Vry148Vw8Eqz24aF5w0cgMUIDeS2lU6cmMhyAAVMk7IdoFpIUk
BvodR9Y/esB1sQP7P5i1z2IF1JLRdnjpuMY44V/SmKdu9R7eMFlil+u8VxRHsamQ31oMGteg4p3V
NSraXet2ZiijES077mhdiR758rnvCykjHigBpznBCZ/o6hePBPyPDOWv3VMoNyKkBys9xEN81gyM
Zb/ChqHV6U9uiR9dpGVl9YPvNXARs0O/wb/98FK51Vlh2KRy/Xh5czSDItuGVQ9NFwzK/zleL1vD
W1h9yVmTFZ1SpSGxfSN5jLaW95UkNzoYHu8DD89yvo+faEJih7qtCw5z8UPhp867aWFIlgvnuoyN
5Vs/FQjrn+mfQNvdko/9PiRqfgHYTyhjkXLAx5veHBIhz/Sq1Ve6XJemu0DsXwZ7VQb8LFY/PSiH
8uJHFeo4/iJuHhj768VsmR8KffIx8cwJaRqZF85kapdvk3JuKAgV8aXzD4tkJCwNa3KP+aSqIwAV
UVyn/67MXWHYqVSfq9zLf0ZaaK+pBcqtLIwtS7SPLA15GzYv4ZHT/Rwae7Kv0nf+xxAFqd0l8zz6
52dv7/razlLHIoxGxQKU5JY+yI0tjCER2EQyaEMzjumYmsuSi5m3YrlaNaLvkhUxA01T1Gz0Ad0v
8nfjobsWnnkvMA+TxSs0fkH6fsMSo2vPaTTV8/seMlq4pGvP0hNhQ36p/NbWSSpltFyHGsGA21fA
m4no9KJKM+753Rd2g4anNTG/3pfkttlEzr3A9DnMDey+2JhR7GDK/e3AUhIj+BvGo9MgCUfIk204
60qm9tqoHUA/qjLOawD6s7gq9dX1MAOVgSaIRqGzPhVS55vq37eVtNp0oXDzb8Zd192Tjalhw5e/
k1cR1JAFjXxYWWzqFvSgITil14EaW5RCW4wd9RwG3/T7EUipA+0KAwlTutES7NLH1/7gF2GJp6fs
05HlOHLSydfIspptXMlL4lar4yDUKTsx8dVFyonijt5EFZg0PRMmiyLVjgphYS4mEV0iNfKCmvOW
gXDaaPXSawqQQGXaWRyiIuACZhaeiL1G7HhIZ+egFdJ0UvKUMjncw94bHubGXZEMzV92dzTRGCTF
KxviO7gOCUf1kktvmTWKUG7TFwS5DDJzg9wfu3OdCNwqZAl4d0aI1gCng1oAL5yWC14DqAW9eX1Z
E/fcQurmOj5pYfQQxvbQq+EYr1viRrXdkjpXC7YzUvHzErN2h7qTqpAa97IepoNTWTEtc6ddCtlJ
Gr4wiCO7f4d8NzKAbQpVwdGZyTaJJZPEZISAFrTeEgz9FUGRNpVfPlIOxscAfWHmvSPw6qO9EGR4
J5yicG5mQBBpyg2V0rMVDA55j2nX3HdJgRgmJgltg37PAAFIGoZOqkmxNsQ9lF6lQym+r07JGx15
L13o2wiogFsLe5VObfnZucWhKUfQuVKQpvFvhApNK3/TiryGVJLiPnWr8h+MZA1X1a6jlLaoecUb
aJx78lW9xTHNDbc3fsLZ6xB84UgOmw2dChrqs5rwC8kNPLNeTf2KI3fQf9taQ0uDZsqVOuOpKCik
aSrOCUriAHJ1zeC+qIDFpfqt99BPlKlcYCHaDIt38UJhdjweq9dnul6yOvGCy42nNVssWb1Lc3Qr
gfXJ3BLu2SmJG2lzlx5u7FVfDTQdOUnXQiSJV3haHbuRYHr0Wp8RB5rOYaOok3ulpOEa055H18pr
7xtGjFEM1Xba9BvldnafMZd2vuVHlzpGiq9dTmLI6CkwI679SNfQ2L4t+hzUHghROhNuwS7oGp0T
dIbFO34lBzpoadJfzVu5Dzz7XoV9FxAtT4UYgNBPn0xaeftVGkjrm6/MGpblhDY0uDjLtn9xmbyP
0BwbrMyWSsDjjxaSQWGOam5iRFpYgtHVr3JvdHHrUMjowwHwww7PIFNNk0n/ZXrc3rIXfbzQLJJo
mnnt+CKFPp0WC70VTOQmJxYowkSnNwdqP67ko60r/PoB5/30TV98dzrdgdPQuRF6lk6UKzKlR4bn
ULSLJNfFVZOeviqy78/Hc2jX8J4GoHKL+h8NP2bkr+iDFojQqIWyhf5Q/R02SHe529sZfRka9+mF
ShfcuHF7tewH4TuSrKLd/CmmyI3LLdEoMzZEtKLi790CXFBwCpt3Var1fBDTrmnyQ24nTrF2O+KL
aZH/heMuhjYUgOVAox4kWBKHNQQyEQWITIMeJX2kbroQ7Q8+Otwji+pX5pHNeFxrz7F5qI8cQeMh
nEw6cj4RS1QKHbMVMepW1cNIn0qf8IcviJdSvfb5ogfT/hfAVCJ0yA6iap0wvSNfNGVZ3TC6gCq4
MXb/HrmnHU7pr8yZUUIW64UaXKwIInd2L8TcZ7Np0o4R+6U7M7+BBR3lWLVu4eReHGKiTMTMfuRY
LNMxgi8P1KrNXUJwftyNgbgrE0EIyRxL5V/hS4wVKdgMTvap5dPwbgcgvmPB3iQ7UoJW6R251SS4
12S25qo/kCaaeQOizK90O5zEaKbLrSFS1SAqJu9ymBUoh9k0drdAdzivHrkOYO0I5EcIL6YvEe1I
luH/eVE063UO+D9ektsGUDPPiyjnWuOAOoxsM3ynG0PsE0I7NHmTPSFiAbWKAjsZ+6Ex8S/KZ4Ms
a6jC28nHlYha0tq12kTuHWWGiE0axcoJ3s4CjvR11Qmvy72Z1lL7xbCAehyco8jUsmqE0cs2xazU
J7omGIjxmepeHb7lYAa3f360gvhaDZlBOS8ILv8CjIuczOh2i8ALVwyqCrn5ZWf5iiZ3k1VOYTQh
pDn4vAe+WLlE1GWrL3OF+l7Dw8tI/n8jCbVs9aM5MQ0/vWw3r4gTencepFNxbtWAnAeuTOGtgWIS
ySrZXr6bZrFo/eTX7AuNZr8QafiQjwBxiAuq+Qn3yty4VG+TH3mBbID67ZNd2ASpFBYY/ftbALH1
jJSGdBVSCdvu0R7VZ+Kw3rMJbzVWmovwkN7YGG3AXdEUa0o7pcwyN56nUELrqKVOTKLJA1XtYic2
TiCPR2snNbKTmLtg3l7vupQ8xVnhiapljIl8s6kkVtTSK5hv1rX5YxAmXz6Fze5ZjODrBydQkUO/
de+KTn0JsgnGqSx0rXj0vEiAJkmme7lMva7OyzhH40okUPjYFfGTunfQg9PU+cmWT87eYQFdbS3j
mIkqqKhm1Hy7CatZC06kLxcCfCF1A+hFoN7+kFpuvg4zM3nubsE6b4gQ4zhHvVOJo/mw8tRLV4cZ
XHOElLiQ7/e/mInIqm6j7FZzH8dx/emQJG2iYeDdmp/P3q6KFWVmKrff5ADGdCrbGMxcet+/MhrY
iNgKUZ6e/7aHnCFyi4N0V7APQ01cYc4uArNe+md3dPVscRMyTiTgk51pagbwcUs4opCqAEOob3Mi
bDZ8ZtJQOh7qqVWps1vjShGdgLQ0mosgCPhvmjME2xtxX8o1Dz2obxS8xuDTFaBQHgKOBIYLNuBd
QGMntTIoFQPUmtoCJpf5zsQ4BTDpNfjMGbiu/T+MdiDGA5S9Ur429Wv7ZeRYGq9HaKIwqqju5r0y
IFbxg/2Bxj109oMVCBrn3UgQryoYxx3aFNYyBPaJQozinqiHj3UEu668PTZsQgWV6LsQ76lqNp7S
SqQzkaHEutRjfrYUtqVm0kV711IdR2XoDslWHr3aIlgsHfzgr/LaqaDmV9+wRUGFzrPY4MTKsYZ8
aomzbKkiBWduKQw6rbFD66xwK25YvUzuYF4Qog+mfqJZaQuGLHDRkiwIiAIJmH2d9ZdGwtsYZj/w
MQti5YaOna9JhSl02w2umoDqpp9lmyRANlTHa4pBymR+8GlM+9i6xwPo/gDWuR4nbjkFr2JXpL6N
9q4il2c6oE4iO3ckdBKiet36dUpMYcriExCyBHHv5trWrnBLp5830qlyXbsPDxyUruokId4LEG4L
XNkytdCTYy1dz7HJ+Vs4F+Zhk7cAXFLBYtlHV8vJ5RuI6w9kS/Zz3iinA65a0rhCbd61XgrvaXVa
Vh+qBcqdjEX6/hJA70OLECl00ngi0TdKIrjmxlMJqAq3H5iVnPSszoRWS5bjdpABcuhHH+3lsF8q
4dyuB4CFwapoPF6A8Oc3c8NPlct2KXUOrue76cAxaAu9Q93Znnd81KDlj21FicjylNeumlXikYTE
jWB40S7HkMVA9ZWFgHsgoFX41FAK6y4OxCfJXIT/RIfQyLW/AwjRml+tPRVDmSOahOurJpWMCXt2
jCykBU97YCZC/BkyRN58R9uLvwKIJU2frNCdrCeA9rG4pGJEsWrk/DuURaaJfDtueyZoULKF7cN/
YozHuLL0s8rNG5udyBHHL4OTBpCHcgXvHIdDWGGr8cadPMk99yF6CQO8aKe2U1iXPl70G+ucf/Cg
C9EWki00AVa+FWb8U4PQF1ox2f5mVKZF6QXEguNj1X6NSw2cBgd+ChVy0V4o3T8CrWGDUOjFw3i6
4xGS9wH0+3xISzhErnMAq7yia7MgMl93/KPUV4x3FJlpAyr3OXyBTFksYvN3gumWg1GdFVScKKcn
xpEpCpq36sVVOUqWx9goZpEq+RGN+CWEjKEWv6/WEj2EMELwfgyAKyaIdyU+UsBScW/n8uwRc8U3
tRAfxUbb/W7sR+K9vZrlxBxhkdGvytWWhmHUE8AcB/xxPWiiiskMy9I3EMhGACV7ILQiFVB/w4e2
Fufb+mbUcvrce1kzJdO0evib6Q9Ny/CaJjzHTb9UTdVWcUlijhVe4V57dAknnGiDPWcS2Sm5+/ZH
9CQqdXeYbXhnLK1roM1uHnj1XMPh0e31jLdIZXZTOPKyvlCRRJ3yg4W0gdGFiws+cP+sIWL8qIM+
T3PnmeSHuVhox18Jfq3CA0YGQ7uwVmj9ZR5Um2Zrtjp5rvR29JMCCpQAahM+QCsdRX1JFUogZ1dz
oIIHwqPwqbnPZ/lh6uNVKJnV6bXb7TipQlVgsC6F37Njv8EMD+qM5rKwhYn2M4Lk0RBmMnt8aGR2
nVCRPrt45QUlYYxWzFqvwjVVlCj0Dq6PjaZsVBOIqnYFWHz8nhEgHUbolzraaOklNICHzG2HiXZ/
o5W4XR0aH0EaW8YM2p1zcJxAPEs+6ezPEEIt8smnOOve5Bfe2I1IiB0WU3e9wdfuZv/4vv2C1dxS
oOGhmWeEx3xkfkuc3YunNSnr12lsyeAsFSe4LL2m9YB+ONlecxv4yEX2m8ChAIaH04MAW6Y5ajXw
Wq5EELOPU7Emk0l8f+fLYqE5s+HLYoFPH2FoSHUqjH4J2k+NZRIKMlQpXdMdt2Egw6PF4rekO8VR
nH6U2bPqQTkAaGEjZJdU91uEB8fPO4hRPNRY48Bs8OxCU8jfWiQVJVXgarHu/DViWNibgz9VLTcq
QE/MhtEqf4OO9rI5jKJsIqDj+c8hg7zyCto7ILnjQApx9/DhcfO15y3RTjAAxJEfTS6rRsxsIVqG
SWmxEuLsAZxMSJJ3ZyvK0ioGm+vrQJNVxnex0WSgbvAsjul790icpBVrSZBnTUYOLNPwaxs2o+xB
1RDwN2FRkkIAIa3FwPgVd7UZPOz/iJOEfaEWYleBekcrYidaL4tw0BzytskKWnetYg98ltUcm3Yg
jvpGLOcvXgGz56Zgvyf1bgsqZQFqXwXCUDeLqSX6eZNMbBNsmDceJzhI192QNMKo/UrAq0w2raDh
HZpr/xO5bCOh7qU0hJ748Sjo649DA7HHTPVKbZY4yoM6Tv0b5nSceMRz5C2OeKGzgmWIskGB/+n8
+VR7lBHbsdsOakEziH+/zXLz/YWE2jlGDmIzQqsD2teNX361pBPJbNV3j5EDcw2YvbOVIw5FymmH
tg9kQPjwi/7dv4Otkz92TdSerC4c3MAU4yGduB/eoP5Q9pCK/RXQ+lGeTCxz96GcwYo0WF7QBAD4
eplfpnkHvMwoPXZZ+WPLHpYTnwYeVUBN5+T1YLeDCkb7mV+i120Au33FQcaIGUPpm/seYP4uniu9
C6pv9OdpiPnTZCw4SXl5UQZ+2BaHcR/KFg4M6ub6z6x7Km5h+v8B1JiPdWRgmem/9j9/c1sSXHVJ
3B1ynZ+HSfxfUSSUS/mg7VD2YefGMnKVMhiEXs0coZ7Y0mooWEXpVYlDMrEOkW45nrQpIJNl+VC7
HvNTkhYGu9pq4S/jlN+npTCmmtLswFzTyPtZt6RPqO5FbW5CYXoKENX4EIgTBwTNj2kEumh/Hc5w
Ztcft33qHeA5hsc5W5A+0PSskEd/FQj0pjupYSP825xuIxf6JPkSmHPFnD2ADSyqEztiHs1ZqV75
CNQbga37XhKzgba/XJIw8kAdHTPtF3kxS0zhtqI+gMkwWSvfy9T3lbg/9Cxww6fdcB+2ETBqI3S8
6twV1cS3A6no6YZ1okEit5se1A+YKm65BGQE6IGP04l2x2sh4fD48JWDO896xXxsaNrjJCCIftVx
Iwo2PST/tW80Iv/cKmD6N5GWnErvlIzzmCZfZwuFdr99RYXphrIPxFJH99/xaOR9srsvM1975175
KJvolgrN5R1yN4NSsENyS2anVS8Q/LNMxgLQmBbGLZYhJygCfNisG6IuukM6/xuDOzk3mvmdVMy+
q3gM01p5BDTY9xYb538U2x89i1uqsuqTL/DtpbOkuwqvfLWchBJ9FxcgcECbjUkEnEfy4CEr8Zaw
VisXvkSeeSl8t5gv0pDOChPm0ksjnl+kq6k7HEmVY/crfz7H0uvu0HSU+T311UkItmPGjZ/b7rTR
88yDxAeu+rwtO4zM3a0zSRDcleaST6pWHGNelBayxLRAxq4ZITJDDqkTvEDQiVVQYM4fz7YQOD+V
JuloFVuulBaMrAGRTWTOaOkQal060Iw/iXirP6aHicSV8tkgdazLcZeOMCJcGAKXQmE4tvctUcpm
TlF6X88lD7w00m7HmHR/E8V9xQ9dbU3RWlcTkqYdKmP1eNE3a9BoiKwQ5zVojYG3ie0HZXXxMzvm
pppAKTezRg+g9cUdr++saxYSsPchskFdkycstxTeNYXSm4hy3VC0BRJujfna1nx7WNvS2FMcNVpG
gRFJLxz5yTLpUYzulmHMji/WqBHshUXykVnzbovqZLJ5eXfDqw5Mh8wJ2d+tDjuBs3XlwT9iSBYJ
lddOmDb/zEWsXirYBOFHHtZh3n05zRqNZZUT7jZw8JLQRnXXYAIrZXqJamsfKa4xJlXYf6NVF7iY
DcDqFV4KcMR8rDJfyEWB1GQKKy6qPK2jvg/29SzscRPtwcpexV8TAvZONxPUc3aBdbTsPVHbGJ3I
pfTfqxIbfjLrhJJUCdWduHvYBGBvhszFe8MfNRWhvUO2vabjd/LLFbOhDCFskQl551madKpIDWpC
UseTd7vb1ISucH2SIG7VD7jxIMVy0n2/gQc6+6rfyu4apaaSrAYHeblztBDAo34o3W1aHyk6CNew
jsc7QafTEIgjdHpZSIuSGJska732R5a6BHfUuQQ9Sfx38EklnF23vO1Vd3KVTshNdJmHF12BuyCn
Ry3U+AQ3UjnBcYAFt3er9BmQqgPckFpZLNTqoZT/wx2vIq9/tuE9pnkzaPklcPipmdEAV29b2Wza
bzBInMjJzIEviCq+tDSniB2EtPKDTrWx12AXqxEjKfNxAKeyalqt8idK/O8Os02vKUTFuwdznAAd
ecU80Vzfj3BuznPq1VbYRo3YNphLIEWsThGHGVDblMPaHfHJK01xc1VnlaGdKv/m3iW37byg9/7E
vrk38PqzEYWUv4HXRbn7fLaBjOHmHNGiHeCWeDzkoLhpUOXKCBTqwYmSKN1QeuBO2/RRid7K/zRW
AcfYcJO+AjHeO0vujJHGYuK31zok7Ig2/uTcB9XxblFOONMmiDdar2UfLMS5cvIHJvyyc//pN0gA
7MRHqnDaukzIZ9lblp1+pDxHvBZSCY0r6pXgnj+pxmjZsqEyOzr41PxBy48aPxeJOwZeNIFtCSq3
fYbznzlRLlFXGzvh2e+igFzbOiONB83VH0g/I2FpSBX8Gb/CcoMSLckC0xgQ/FQ98L72zFXJPm4G
fD3g8GI6oN3C7vl5f2HpGJgDd+5rHXV6IXyqAuuj7iIown/JjtfAxR4suk9oVqjs9uyi+5nvRUQ3
eomMFtG7eetQEZUTd+o2unwbMaWGJgM7G1KrCPj6ywJlCc2snNUb/bo8ZKF9WYVN1xhX7z1ptI63
9NzWXjxxJcALZYEO31ps6q0g4GjVQgVPkaVjxf/EQEZeBhBDkaOygBcNI8SJZxD+Qk4UaBxjo00R
jLBdVB4EHwW56Tzk3KSCQ91jOiOHeKRu9WP+Tn4a5+RZKIdjd/Vm7PQoLH31bI9TtWbPijowqKKU
po5rxo//PW+MRmI3AAdYoS99u+T29bNF/isNQ7HEpMpijbT3c9bQ8L3PB8hjwhgtLRKDORoKSoEo
4ID6GEHELA39gUsTbbQU53hJGr4384WNHmd3gH443A1+NdG3dKyvndV5YnbjDmkaYeCzVr6VJ4VV
JTWZNTZhjkn5hGcC/P237foP58/u+ahSHTdBQN8ibBEjhlK+t3sifV+YywuIWf1ExBnWN2CJPvfd
dCnFrf8PC5FOma8gf23XRDW/T9oxjPDl5yYq/nXkcUG5lfE6cT9Hp3HfcHbpCVwstI/2Uo+WVQ1S
HBUH79036pvey7sDUvjS9F3mwqqq2S8ySQfNOf2x0sBwqnOeT6pGMnYYuUpQDRabTIbbhunoQ28G
d8ozXdA/hszRGL3R5sXcba72rY4uUB3LRedeExK2xvCaLSGaBrcljAIPR1y9pn6pHsnaUk5ICUpz
yB4OhpGeyAfKlDa1YsXn7F3bXCfVHw2hZWbiRncs0YeY509j9uqXWe7t7Bfe/Ncyn+0KQ/wVy+74
p2qaUXOm5aeFbwPYEaSFFzTBSXRRRe3P2upjA+8LijqeGFqpYTErQq5q3AsTDTye+IPWS6qY65hJ
m2Q9pcyCavTTcLW7okWiaTw6TwB1ufaxMZ24PQ8BTj3ergs9d9vzU04/Hen42MpivP8GHb5cyfDm
1Pb27PiMMcoS8dkMr9L7akPDNpcMbwRGnQtrKFis79U128ne2ZOG3soDTumjVNTv7iHucp+SrceQ
vclf4ASw6Z9WMZt4x7KeyREpth9HSNnYpVe5RD9OMEYA7Qlao36AglsIIsh8RSXHZS1VTkX/X/Kw
wIfSyd1U3OWPuYNf2r5V9aWwWiclMMcc9BbQQIYvFeGTERO07XXxvd5DUh/e7/eCDJsVQMXYoqLC
B1G53zuRAPwFGMyadUsBlr6tmWVCY7vHO+eWBDKwbaXs1l3YS/kpgptCb8z7fE4UeVnLj27wxOIw
MH64D26nEqe3KmZaKHPFgQvb8Wpw03P4vw4yZYPv4txY3/aoq4LVmO04ncGK0pTb6gdx+MJAFOt0
a+RAybHJVKfH6VTQqFJu95wK8LNzGbs1fIfROa2cLh+aME+IburlE6sG9TJ7tlCsX5hbj6HEmXKg
ytDWQUgXkoeITdv0XDGEYKuGhBEiPGcXimODOKM12UM4CZ1aFuv3AfK/hmc+h7uiVyedzCKHR1LA
cUUqvL2cjFJ9PW06B6ej1uKXxcUndBU+3S/M2BfaUhV4D8Ya9dXgdgN07v906Ox698lZX1n4OhX2
OL+rqsZ8ipEzWH8AVD4ySX77OqDcB0Zw0oLeghtDd7jKSve43jyUnlzI4ckGTeZRHfwPm6YrulTI
PAE9vPtZoD6QUPKpzA2NjDbEQnakAz1QsfXTKvgzkC4CpuZuyMjJFWyQw1jUw4paJRFI3ZXVYN5Z
2G5y8Iw2fR/JxWYvCGYVPhYtViN/uTD1XUTmWtHqmhruNCAzB5YQO4xpI5gnxLJ+zptBAL4cSqHr
7XhprpxuxkTL3bDqMjZciP0FpkhsRJ5DglbxzU2l0Zacj4Jd0u6mBdT2UPRAu6NjJwdqS1HXah7E
I0qb+ex8w809sRKaTlHt9gh16JrJT8Jd8G7r/kH1ku4mW74vck31hgEEaBnyhv525tmaHZsEDlDQ
2u/UGig+3zqiT/OtMsAXI9WoKdJDuxa2fVUsTMjk8Q2N3g45rvWkNsBfkRqpELX3HE8hrMuNEQsl
F3Mbn3qbfo6Xf/ET2gQAmQdfMIY1SCAIChnEqQ110UzSeHaB1VSi/BlPgUnEyduqgVs6ASUmUOty
G1KVp+WDGU1GRLM239lRxwuBtWAMMLaC87BHTKrfc8Qvyf22O/fEavOpVD07qIH1xtDnNPe1qSy/
ivqUK/PQTJU7tR32WKYkbd4YNtAIhENuSdW4UpvhBr1Yj1YNbVH08UdwzBtZm8NbKrbUAl/VcZih
lcTwItQ8tpu7jzRKuUZkwe3uSNMqDz1NCwf6caSc+C3507Nud/1whEdY+O3hZO2+KfGSV2QsUCaB
r7X6PZDDkXtJa2/g/ep0EvTGjOj7vIYAAc2KiDNhF/ZstCbPg1R6EUC7u0gnJuHIlaSD9VMDzBiJ
fmmQ7a8WNpNWGi2rNhWXgwB3F28EyEINw8PWsfGBkl+vicThMAA6EDLgBBO55ZclmIszF+wKSkSM
1wbyv49BCeKY9qYxvTvRsRDSSTLLoU6GSJvurCLisUuOZy6ZQleP/BEIUzlRjFaFDT7/tSnK+cFx
pTlGNf4J5uF6p/iym31XohoIYIlExyCgLsFmq/EqkrOrbWUCTsVzWQ6PLSA1lnn0AB12ec38f6gJ
AYS1kjJhniNcNOGJZv15fyh290JGdG6piVOuwXZRobvBZ5o4MaVxntT9UC8Rv+5T/WbH+q3lHu1I
6MQ4ChAk3kARi/zoMXtSvCzt8n8zlrUXSWqAfHMWjNkPlHx/qBwIXywwVBgnjVnFACGMTcPyGzbd
dBoHdzOe4cbxtNvYIMIQPSMi5JOThpuML5zjyMz1tVLUXEwj2H5g7mvolmND8bpeDt3Lcc3k/TjL
I4zKMMLFcjYxigkvllz+6PVa/dhXVPPGrWV+91Nbzx9MB90wNDElWq9ogM3m2MY70nKX30GSci1N
ZWBS68QXUxgRZ1JNHr9k0Ai7WGuDfg3H+qinnf623DACYqS09VJ+6hD31DmiwC3kmahcp/gAFpmO
OKsyzN1KCuOKvRj2Hkzx8CqV3k3J6Dn4JIusX5digHmkLp5rqIy6jqVEXB2ybgnOm1ycDbjGd/H+
0cdl6h7pc11DHtAZ698Q3WS/05Fb07coYj/zBlwpyTEk3KgUcxUMs1S27I1zNJC7/zTZb1bCt9H1
K7juyjP5Y19SuVmE6yXxX+DUU9kpOPiJemiYl7S3aqp4BPTAAgbCO8H8qq7jympTeP960ihN6iNy
32dyxwa9nFDLNDLRQE2mu3iiPZR3glmXPw/7n+Qc1F4VH4cqKOU7/Zggd8anqIeIVJRvzyxXwhrL
o9n5N0qmM6OmSsLQyHo0uAQmEsUo33G12GuBG+gbaVWFxv71d32xdGXWB0G/jzPf9LK5SE1EtNNH
0tbGwRCwtNxpy23Yt5pM6K0QHVuq6TDX3XiqtlVU0QGcOuZoY2cPDOSbwWclLhyifHFoUYAZuNzn
IviBUIMdV9ty2Uj0N0NEauem6s5MfqU9bewbv7l8VMF/rbDi9wSFeSpQiDGYRoaYZkoqu5ohikCf
vnwljBdJU7Nx9rJA+uQc6NfRzuVK5ZFZ+ZPhzOzeFvWbYconJ3uujzG3R++GPpVaCiif7ELD+xHN
tyI+OKxbcav5BIVerXS3w4eJJM3+O9JOTZ/yWH2lxDicMKPHfW8VmrAPoOIkG5KtGeVHEwquYbzV
JO1Caj0mTF2l779hlXYKSYDPgDnDXrCTt/fkMdxqaG46QZ17CSG1dhoj2JwNjOXexQuyUlE2k0Jj
+bvuU8DmhlenxGEnjarFG20jyuuASy2/brt5OIl4ZfK2j3s1miFBVRg/xcXoU98J04ZGAEjr34lD
+57an9IVdZyNQ1EDc2WQV87a4Pqc808pGUSw5jWm16DscHUaNbByulcxiyhCkdxh249ZZ1OT9GZW
6aZd3FrYDjcxBWEEjtIzR76zN3kCJ9EyHg0NHk9pYb7H9HGAW+CUdZ6WtxMUfSrhMyF4VbmHN4YA
F6OeLh5f0Qg1JSiOlG0HbN5RIi1wsw1HaKmIEIrEtz52lpwGMqysmISaWlClWokshvKc50WxZBgj
kscR9yz8rY3/i1Fsi7zA+SML9XoWdSzkcR/bZox6I/r4RkxeTaDuHGjGHIbHUxLkQkPqdT9DAXNm
91yHi96Ut6bghIq9EKpP7En1DbhbYmJK/QaLmd6V1fGkhkI9WyI55TVLmmtAEEMWhR/0Se7fGt+w
BkiBUQEbK+lVUU1K377V+dgcEhiYp/yEG+w8xfhIbNFFieO9YbG6PrJSKG8R8nohdY4KqRy2Zhub
e+sD4hwJ30R+eqQCSq3GfmGbSaPs4zXKvKhVeyGyY0topm6NnIHujNsjPfxHWklLKoL7NIywIyOk
zxzudR0IUdIgHkGEYymKtzwCGCVJMoEkkAk7j0lONmAkT5HunwggLqUoEhVmm7xL/gV7MZKdLFEL
sp6yk63w+Vg1+rUO5HKRzwVmTJAuoAolpHqCOG6H9Hotxo1IaElkVt39fMV/X2/GPUbme33ueuMT
An9mEaazaju1j+U47PzQFA50AhB1uh5/QEcQ1pTD3+5z45kh0Hvo3QhsnLWeGVSJtvmjNzGsID6N
F8mJttvqm81fPK5YqA/KQX6deUs84nA80eNxOWB9uSNp+77BFGFzWf/OaLLcmvU01CPif4ew0fAa
Aj0H38vrdXbqqXeovdC40YIRIln9HjzSAq83l6ixwI92gx/iZhlcnrAINpF9IwqCUer05l3ytDpE
ecFGPu4fTCNHItrOdt4vddUv+fTvMjR3PBUy/8omy6V+CdbeJ0u40OF5UAn9EVnQa5H8ObyNkCG0
IKZ7IhY4QrxGwHvJ4ZlSCZtaA0gjatH4gQQQd3RSEW9KLgnJOALcJob06kOZrGLjL+sTk0PS7HMr
zL3MA3JRzfe2yOQbqWMdBKsvyZGGt0BZ472f/EZuC4n91BCt190vzE0TE9c+kFXu2VRMQgCBQX7R
txkP8sqS+IhKwj8oCTF265GKl2E9+uuEXCqbXZSHw5hSsibxjSEScB2XgwlPahlHk1J1aqmbClss
4Kzv1w8noIo9C3wC1UyGGhgBx8yuHm4OymSfkcNshq+oOOoIHsOI7gtPsRkGYIUbPS+O3T46uYA3
wCUMu8AcG7LjLGSN9/3wjW/4MK0JC7giBeK09FTMAkv1qmyyH3zJNGO3OTKpWX3gOH8RNNwin2Dd
VBkA+NMSOhqmoebP2vn43rjBDTEZGcS++IR9jEa5ydpcbG4C5ohAR0swzXWARJJhT1N2OOYmBWFP
IFS0MPIH3QzD4ABXqXixYGXhHsUgVIP8uPQLqupYnSRK/Xq4/u2vUTkk0FkaEaTHUNYNjILxCpjJ
EHqrWKCNCHrM4uUsoCUvD2Nb61A5OEw701PR8kuz+b3ZnSfyhDgQlE1s6VgTy6qGABI7l1gG0BC9
hFsUrFKAc2YQy8s3Zve9yID0kNOTKxanBi5yToNAmgwugBUWAPK4h2WIjs4/6AMYlJ7afmeRYcNg
h6SeAwatCY+p+PfCdi4ommaVWFQ+WEwacHFsqIldqIFvj5low4oXDvr7VHqhIewwdMrzCmJbIdcD
ML307IPTj1NofFpjfQDrAc2A+IHR09e1Z6oEeFPifr6RzSGWt4fypT954ANRKAPbBo2nmbCwQptv
ewWi/l+P3kSxK0mfDZkmOZHp+RZgvDbvfDAG8bkiiIbKde0kmv0u9Rfl3jcp/oeHzuLxUFHQ4Q5e
sydnNz2MsFU/DoDxnVRvq31Xkrz39tn6yU25kLd/zt86lLc2u7jfN348B25AdZrIjZ8Q0xPNUaid
u001MDqT20S15IFeKTEardUjU9mfygot20DaiwMaFRbwkwXGyAz99sJYqeUHLL44idQm9kLAnVpd
3qLvsOaF0f3Xcl/Zz48y+DKE86+rZFQ32S2T2NYq11hU5DwkZ8YvFLfFIaBgTG5XWOHzmEK0VzlD
r7bPIP15OACb6DNGjIszZXESqyDIDuNI5xipE/uwj9rEFTn+DRdADlIodMi81jw3b1WLATBFyQix
qxHgBrVhKl++o3tyXw/7MhtVk27zFx0IO08apyKrrNC1LWQgyzEcMdIUzmKRyfj4zIbYI0Z+2eYI
UgVu0WjflDj6561WZ1MG6BsBZj4mmFTwNAGbXKCxR9dck1rW5bjamlZn0PKHyfKxP/hkcWSNc1Pt
otInCdmeMncGkvpZ8yEW/NmiCDDbEMFy5OeSchn6E77b3leOC20Kkqta/+dkeiDo/GGHNiLiZn25
EGv8pYoWJTvmSVbjoZ4Y4SKhDf0Ff1jsPQiXFVBFLXat8nr0sBZ6yQaGjOFxy6e0sxHY0QI3io6q
pmJto2cu2/beZ1gTNJZG9zSVuleOGBaSIcByNNPI66K68uKjopWO5gK1UmGSa+BYau+Fy8xn8w0+
VYRwawBconqDClD99O2ixceRhBxXH2QrZx089laRiioh9pnG+RoN0x4dw1S98BqUXwWGz8BD6oZ4
r7pP7C6YrAU6WwYjjo3LHsA3t/OshoWT20mahjBzbmAlHT1pM29pXbc2t7sIzI6oeYC0jNTEcgZK
sn1liaIJCK2sRbuYAqXaeI7Aev5xEENRe2i8BVbHYV4nXX7Tx/tLJ2DHBBxYZqVVED/4fclb8WMZ
rLpQYNvzmK/vBSaYp1A76xDlYVzsDPsKcPYNBcUmm8UMzVcGl3R0mxvVg5mJxvQ5yvtvibN1jlsT
87WntvRK1/fdh8H1aPbEwzOLZSjypmFwDe/+WlFG+oqZVaoTpPN7dKHjkgjgWCsAd2Mpk1DYIkhT
R/Cb8ppvajJjQW1Z3jWQNlIMUiF8TJIDW7yjZ9nARF2YiirUvJ9DtRDuQIsEMebkoZ8HzLekT077
+wPBG0JV09FLaGVhkZW0YLHo9HKsaIRyFkDPrDVjFPdflOdilFB0nMVMc6YD8K1Q2O7UQFzsSCrN
IXhjM4p83Xpo99YwGj6XwJpDYVkKnKVK/7B491R4lct1z2V3apDLH0tEFBthhcGbclXQIG40u8vx
lA7kCR8gN3Hjco3MogETB7xUgse5IKyugvLEUfU2/Uz5q/nD/Ai+XDwKHAzm6IK2mEMf9MIcokv2
z6sejX7sIY0cONdzUr9vN8gUInzEEfiTmajkdi/mEa+tp//cgwvFkn49XAPVFDvqpLAkBvb68PU1
oAvBU+kndcA9XqM8nFFLzQBlHw0GswQMVsQzFF4iTNnNlYJlJ6hYIdEFDycS1PabuJaHxnNsrbru
MoI/l5Wd/b54QveeTH18RzMG0zIjS/hZaeHanLxOENN0e11wD3euywPLeuc9E6vZowp6BM1/Qj2V
TZUKqNh2qlaZIZHZ8nXe9KEMazm9PGK2iGwvl5J6MFZUtEjteh9r724F4IoFlw9bdxDGMV7daQl1
v6Et3MRhMkUVC5exoV1wc4uETNkrRkcLy44NvvJNeJWeoWMgtTzAg7LBXAnKA5Rzds7HrpJ0nYSE
73roMOvZCuP7LCdbF4Ci8eSuf2SttVZVR0vlTb+ZcUwQ7474lnFiEKmwYhSx8ApQUaksi5v+9cp1
/8DqkKRjMC7t1j4UhIaOkPwiVwEsMLKq5ji7LA7/NFATlWFTRX7HVxlFDWI0Jp+rp2PIXWr6Ris4
j5PHFe+aqlIMDKHRnoYlYAwalpZrCMzYp0JsUauHRx+B/c7sHptxZBL03cxwayrCD6YdhmHj4Rhv
Ch1aW/WONhoM9G08z+zaxky+PVKW0UQiDz/nNrZRJ6GETMYxmQIWwt55T+UW/1A3xqm2aYPc0DCP
ioQDLboDsrf9alupn68Cmdm8fxq4A8UAoXWLa+8ExI1KmI4V2JTNEb6o36szjQaQrSf4X+KkMlt+
4Z7kvl/lluhoKq+bny8/tR52mPmuEjwuKOJiJMguH4x6u4b6FWVqYkeX2owItLHh4qV5FMyf23zC
B8Ad8F6IBT0peqP5lFcy0ua9OIDcUyPMYu13Ld/xKd4xQMnngAti5SVj8flOlRGonBw+qSgVx9qj
GkEnKa+eFHNCMj0SPYLsIMtERE4N0LYQDLscsv5CcnRiTL4ybIhqLp9QxtfbUaTSEQbeRXg3+KMB
wSxJhETz5v/CCukHA//CbwD0n/BhYEVzZYJ4prcGBapzJl/ttD0x/s++uJZXuVd5PGHazqrRRX3D
IRp5AAl1dKIQOXWtjK/7+Ib0syZHE4EN2hbte7iMUBEDNeSoaPN1wGobqtfeBA8V7P6snPy+JehN
+Hs19vw44yKFs5n1PjbfoTvUQpcVk3IV13gGjZ9DrR8LKzF/vjMet/FMVDKxVPq5OAr3hp62bEvc
O91scRvujTK5gVCjTKpDenoERWlRCYeIg+yhF3L/FR1o9f97bfJ91y+hkVqi1+EadZmVuGkHE7y1
ACtZ/f4G6ub/5CmrYL7PzV7AismJFWsLgqHFmbtVw2E024+a8hwber4n9ulBzL9XQViYOb1dkSiC
3ldXYDiexPD7wL45neOVziQGIBd7YRS4zsaXBIyDbcCGEfPPp+AnFA/mPkhzLHMK69DmQ6Df/Olc
uS+HTuopIqCtWRssM4EYhIQ26F475oiLWUPXgcbmyXTLiMCqzfM4YWH9ULzp7nIDW+fIzDpRWJN7
ccSTCs2qbUKfnpVGunBDmkSN/G76GdAFowWA4hPRVqu2skiU5M/GL76ISDPQfkGZRj5qn83ghifu
hAhqrFXFt3sRF/N+4JtV1ccq8GhyjNJmGwerpGfHEHbyKB2c9XK1zuvEqDzI+KICNnpd8hZdpMUg
l1KwuKymo59WIhA7EHQwvtUBAA3UNPKU326ZS5dps4Mg6MuBRmFcCTGGvT29OMGyc0JBe0IkO3tZ
Bxt3cP3QNyNDYmZtexbykUWx+f0euof2mb5hrZ+Wt5cEEF8dTJg0I2zfA4xgRsiBdx/y7JH2AOYP
MGD1bnoKCAcNgYFFOjiKtrxvxDHByr0QAnTB7UTZ0LFf5y84XNS8TBIv5rIl/eF2GTmjwZiP61Or
2jE4MzN0WgjJRT9U/j5WSi1NqbExMQ5obbLUW1bw+z78DTMzobK3uBj7VTZbR0eJWKaKynK+lHfZ
ilc4oozTpk5fbC7BZGqqAqflTPCBXUnegltz2cpEIAYyVAOyGUgh6IwDYCpvj75rU0Heh6mHtZLg
ABZ447BpMmIDwv4mzkan5Hwyjrhtu9pLsu/JdT3BZsx4DIcBaH3yx4972AXwOiuKttR0MAQSjJ76
RUrdIAh7jIbgkZvC33ThsXmNJP40FqcbATt1THKbPaRZrnfUdyIfzZ3e/oqJGhIIzVysaEuH6PB7
HvConhFfJnnvYzhrLbaEcb19Q9GCuFLnauvzF2RYH5hX8iHKgN47lWdyKqaX1POMEM6yvfBUqJT9
gHJJxicUmco9BvIj8/eGmznEVgLccKpTAAns/oCU64dIRf7ebPlx5qtIBZOn5aSbgI9M/Kkz+fjG
Qv3QPc06+hXBqT7h2+KaDblnsnsSKOxG2zZBuqtMRm6Gairnb15fNKfxu2EhRU1B1UmVH6UhrA+5
To2zKyxl8oFFWy0Hfq3QTZl6TIG+4f3As9H+RQcHf81sXu+S6cEburkLyW1Z+klU4sEmmy5Hvupq
DX+IrJs8zS1I+lbz4jkW2eURndyharY/83SdGL7P0EefFTGzH/CfjvSrnfUvxaFaso58trH37+tb
uMoJeLNqJ/dhbtESwhY6UetY/MRSL7CINTZyLt0t/KyVg3YibI/crLcAD0Akebse203AWNepyQIk
WzJvkzv76mIg0yZ/7BneOkzoFo482bntFMLuu5/MSYHMmh2lsaSGNSFgjeYLejznMv5iGhefyLnI
iULRII2R6gJsNVuA1py+5NYKLWYG7emZAIedAxUwxND8xAeFYxDdALNafkNKajRS2jzz9XFZTAgG
aiYvmOmgS7L+7X3hUzJzrSMS2NNlarrBbdgSYa3t6JNIhL4FOdnnTcj6SuENnZKbx45S38x/mgLY
SjdYUYwrnIpuGzwqRjBSSHiUu2HDnBoheAK6qV3WN4uylHamXStQJaYtH2WYiJPVgFcVC3lQXsD5
kVnjdhaG78oUMimFbbqwqEtJOj4mEWPYNyRBbCDFG3YUw700te9SUylvyHyk+GH5eRdnIexy4yTr
eAgKEkUOYm4nRM0HQxeFlcChDzdQaaOLR78lV+S+omif3ITBomLdkXLGZhzFsl8+Zcv84MJPBZbT
YTi1sIc73Y1SKvY4jjwPcRdvZxNWUsrFwTkyu4AVhxlImKG3upYT0CfPhIxvdcg9htDEmqdkcVEc
ub1WVdAvGf5QkWTdeB4HvOSRNYjInDGVkJLSYsAcwDmAmIK+ReJC6WnT8G2KDaHDH7ILvGj+GXbz
1jXKe5rj12ot1ab6GZxN5rQA9Mpt6hEslIY+2YVO1yZT315fYDz84VIwL2/wm6aiZjfVokIz/148
pgQqKNsuLKbC+3RMYNYqDaJu+awq4XVBhHtN8Pr52z+kc3ipt7SQV6GDNPC8OMjbiaiLV/IzTWjv
QO8nJ7EwqYjLWBE+oC/HjIkQ1dt2mpudh4zYE+lyutnGouVf6VYlt5TIum9cpMkG8fe7YS7KluMC
UyQ+GXuscjABPuVC/QPfGU2wI9DYjdctRGY+ZGKzdYX40DMx7v+ozzzHjdigP5ggCwz1HHbqb5ev
dts/gJO+LirZ23ONYA5hxoAMlpsPy8cFTD8TZB0ABPA/uV5ejh1YN5bYe3MZJoND8xu8P2421LXy
hchEx24eZ1rb9uMSaATqFedz2Rwr4GxDUOwifCZi72IcqRQEgeu5U9enbQbF7wEY5X0Q/NthuMBH
HahHeWg7EJeojZcLGEMUztDExqJo9nomoxPF0O9jKeImWSXDdzjS/qcb2eHq40qtkoQXlgc8TSoW
DoriuX20Tcx/gRJ4by7C+i76B8eHVRB4JEAPNHIRbzsjPd7P2tahyO9OW0tBL5t4gs6/VM4F6WFz
g04tfQQBMFvVNBMJ20xBZOAFb0AdyC25QpmZ3p8n8jgEoU5ARXtykndQ5xwnFLO5GKdGxwmQIEWf
N2YLMmD1VZCpocmtU43+XMLP557iwD3aA/GTZh2jRg++GXIdlDHyt3a1xKvh+KYa4VD94Qp94aG7
H7K+CD9IRUvUKgqZkOBIEp3eSvQ6IqtEqHEr95fvpmckJfiyuX4nz1ZX/HovtUOe6HSNFwQXC0Ym
ZlRzsWoaSHCnI6li6cxYiPQ/IqS1jqTO0jqcrhhBjT2QCGSkuNVta73/6ZtiK13D0E4I34xD/aqf
Eh2iHZ/8gnyrJoCm/5ljR1kgoun+4RNJmS1q7T3O7jO6vtNeBKLDCgVOJjoWkKVy8s0rLNsZW2tR
nsqwhAMMtc8YxvCqMr5HjxMHe1N24sB2M+LF2AxdWNdSqTtJy7LL69PandOh3selwNcGDEmY2D+7
tLeIn7CQIwUxfEVSX8rM+10Rkz7S/AZScIn8OG4Az68FeMXlPLBPfxSMxlzJxDWM5y9vQ0gMcTSy
HxlWOvznk+JXxLfOyJVVtCK7wfYwKKXZo9lTFgisFkycbPJYZ8/Ous95VnBgbgYxWRiggb/jQISj
TV6f7kx/SldbOwBEVKAB1IMW56tAqTnoLhhAb0miPjXaV+kKxoXTdZCC5GqLzlY24Vk0HmYhVBZz
J56hw9Kw0MyvZsHGHV2IGBEC3P2N3eV5qLOtluWEvsu0JvPleaJNMld0AkrhOSG0rX7hJp7OJYbu
fOROwqSv3n+wQAlkBvTUC78gWyhsZuyianGunIU6AG3DEmBvX1xkoPgBZ4AYsiqN6FE22aDYCKH1
qhu26TficgXry2xVdYruZ6xEQyBxTLxI3tFTxGLRQPdd7Jve/9YIATuHWyiz2FwpYH+tPXR/Qpy/
PjK/DdQLBR+F3qSXJCHCWYFW3KU+HTN6/jQ1xcfAbulRf92p6f+ryxnaLE0KeJvpANtJaQ5P/Bnm
l8qTX+cAyP5ooYjAluERr1SGnG4yb5PmKWWHzeRTt6Zpe1padB+Z9ledRlrDCY2SZtZ2NXxykkEz
fvrJXko64zmRmtk70fX9sD6fvYrjTptZRC0ExFJIOvgmrwI8iYQw/fRXdQYSTIxJyPc8KONLON1F
0sDTbTe8YjqkZYf1N4UwlXQ14hkRVKvx+kH4OjTXuRQSGwMLIQPzufzb3d+0Y7gIRbXw4vdsdnWO
lrKy4qiQD3CmdbdxiO88B9m3KXpM3cdF7Y5LeCBWQIWHjIqm38icPp5PDBXZjiZwazBENvxV14mw
XphV/XFS9Qr/Up8IJU839hpX7S7OloOcx4yIetBYFTT8p2McFq7Zzm3t+MpLwAw2j2dCJlT9uKXH
2X/2JGaEO+YEkxVg87jiClFaN1qPpXIrYQ5oDGhwnQ5SSEICIkoVao3eDyTd0PHUZH7JGd3exIog
pNyrNSHfsL7AoANs+c9Ge0dV1FQk2ARPGzVfOKaDgI+F61nwQRnzpnScd0BQ3DCpU/pykRpxSx6f
WEpAynwHHO2IP4WCAtGTjvebnhfoqSunMmnLm544brrrdNUWL2uJY9v3+RVmwgl/Z3mRM5ejzCaH
a8X4ZLjyTRuU+Ot8DAQgTpuX9U0sb3A8344XpVbFdWS0joaqoigyZwlfNCuxzIzC2TXhk+5HGTrJ
TPnQIK/+7DsUaOZdIcR5SOk5eSp6EuB6Hjd05I4HjnwahGotf98q03CIeCRpYJ2WO1FJfBzFnl3G
luDbGLSxf+TTWnSqrEORMBMTF8NxXcr2dTVZopN2j1wG8h+XaK4JuLDbdlZT2bZnHCI8NaiqKjhQ
eox6fe08V02om7YIGWpxOtdruCfWE1wpVFo5crtyBCsC18zvutj7vHx8IL5aAYAdGYyvo+yYKqaX
5hAktNeFZjVGDgS1z6v0KItmwWRAJA/h6n8C24+Q5znMrVI5H8Jy+/RuANnM2q0X9Zklyzf3wDAv
p2w+5IuO8IRtkH5cSnk664/oFJLfsEJux5dx7hUZzoNkXX1wdHPZXnvgss7fROCk1dsFPgTAlwwg
KGSJVZp/E42w+wQ93BaoRlkCYz+xZKTY6qpflpYowqf6t+ieCgnjPyCK6tKT36EEr2cQziTkOEgI
u/bbFjhwOCBzPFOlb0x4SLJVrO8yw5vjdgf0eu6SW4RjTKf/9atxq/CXvtVbI3VLB7CMPCVBAAzT
UghBL1Q61EqaFjRuXKdFyibHp1cWuiZd+HY7V2Y6nvg/TvXwAR8nsO1Hh6Izu8P8NVSR8S02XqtH
icrABtoAAfbIzcyzxzvLWS5EwEN7NLvKGC1zfL923JgViJoaY84KxpYRezy/Feb6ia+JYQM83U99
6hzJNkfkleFeM0Ux6yUbL7Eg8rDBYAosZWAeCTJVlszJ/Gfg0Z0mQI5uUM3wjK9XuAj9zzmTcTjY
lpTzuclWYeYDvrAGa5IZ3IPd5etcZh4Zu1jqEBzL04c0oyFJB4ugE6tnwR1p4XvWHGdrH27zDdZr
PMx801DWqh2yQA2RKJCHlDde5QxY2MYmB9RAOSORg86GAEAJOYDxj2x7wHFTgeD+oOhecHP56T5Y
PqEAN86YZX74eWOPXgvWd9enb4Nt5+CpV06kZo8IgR08Uh4IDZ0auEJ/14jEthBIMyE2QdNX5jDK
bj5ttfuz/uqAedwtbDyZ6BMQLacjwDAOMRvrRRkw43xpcYXOATH/HXXhToi620VorBxPL4cCbQAB
hscA+oQAkqRN+oRdfVwoeFCQOruMo18TjrW95VFIuhBzAt0Wp5LKFq1plh4Nz4BPnljZ30SAbdov
v+UAYwxNmhZkj7NU9yjgYdjgnP0+EWhnGWonk9DMWu1LAtiogpnnI73yCUORjiZ1DOfVyaD1QNcW
ZlevBtkc6R/XWwLPc3jRG3KVq5tlb3mJT2V6qv+gqEg9GAZPg9YRK36EtZIp31AaAxbgR/BfdVmK
xhpeEFT2nFcMNQYuxnPd7EZ9gZKuu+t7QFjsOF+HnfWNC1vP4LkO0KOcU5uPUsL7mX7mO5QmfhSU
2bHiNY59zB5oMUiWko7mFTv7O/NGufoTnLLR6gWrtIecZhecqQdgMO28/0WICOczKONoc5/VJnp9
17+iN83dhGmqxTPn26EKhOhQ3tmfGrIVHmbwhxufuDPc1sjFRFrcfPWD+4/YyKW70O4vRTTXhoZ0
GkE9FwYYzITzN52KdPz8B6e4U4OaQ9PEG7kzKP07DRle5V84ZrLWHKO9r4fe1l/wBCCjCPwhKPlP
RG8UHQurc8DLbY+oGV1ioLvlczlYx8TTRmVDVDCwGSwq4qc3hHQqNQmdR46MerandiKTwi+TyiKK
jrO5wo1ZoeCT4uz56P2Rp0W/FnCY1uHDvLDf570ZIIE9wpcuP8/k7jO9QoB9cjBiAIPktnKRPyFl
/xBlW3oOqtH6ESx+6BMoKvrXJjW+K9anjAUtHOiAV6WkmXqzGWHc46xYYcVQVd+koo7SjiXBA1yF
awd3YafqPcdbKGJTuZep7kpT1uqRDkRsOh54O6FzjbvuOPLfnW1mCEmqozlNjeJ3sO/4gwD7kR24
IlNZh98P9T+T9qB7fDTN0YFEV+8e15Ar49s/lGbTtDi6IbqyDHsCay//RIMwleHnrtGE+3prC70H
O/c1V9i23YT/JOtg8bgdGxVGQ+yutrzffX0ynF5q19cEnQg8jddWPKwc38yiZIHehPPY9qyYdjJI
U77/qAwPhdMa3ngCeQ1FuzRLfLF2r2hIP5fyM4qqY3kK12VXBrCN9wE21zliR63d7N23gKUmip7S
JoqgKJ7VsMdbtsmnda+h5sj5Tf1w8xDFv/aVefNgMF40N4nZ2anMrAYi9nve7TiokMqivwZ5f5OX
D1oH27UFxqgUrmEpwPtJtGbkZXngGw30Tcm86rHuTith9TvDWW+JS5NQfNQPVXpXchWaoD/ruEgN
rkRtzOZxso80jdvkcOZDsRK5RFFaS2cYX144KNHJk3YhGtRciinlaoRfRRCi2DFo2gcE5l3T2477
hSwR8wAPfdykQ+VMlfeekoIvK5z433OsnLyPUX3O3kpc8uA4YO7YKiHWAXApXDIpoRyT24A3jwz7
KcTxg9Zp22MfW5eah2VAYzuG6cE2RDCAQW/R29jbIWS9DTMSM1n+iVDnoDUWoH/LYn6g9qmL1hfl
vP5I64vlTw7bluVj0xux0agjRWg0PPGCy4mqmUO+E6sW2Q21PjKWvVcaIo4nkP2lixigK06XVrdL
i3sXspZJCdcFX1/yIEIYagDx3LQcrQggLUB4fR80CUBm+RHe2i49eIPtkDPRZsyiY93Ihj41vAAE
BWVYUpMLWXnERMW4BpeoycEUD4wg1KLndf788cRVYMM9L+9vjtrdB3+dWjpopegvjrqjs6Xl3stI
T+JnWm/YUqHbu0z6RLPeAS+zn2W6L/SEmTvRzBYuMafU+4ZNn/eBo2IgM6q2obNERgd9CMW3kXLj
YJCrjdUY4VDYppmatkY6LJVZ3OO1raOtlTewsxZmVQrspJBzHgfChO/yugJjNHR+TlH46//RLygC
wtSyNv63eH8CRzgei6beAGE9QwFE7UADnhGTps6vaLZaEulWbpVD7IatcOVPB17cC18O3vfd3SpG
rHsWf6HO3lhmSxSqgZ4l1n1n4DGCISvhyjCLPyuPzODFzR1oFCWMw1OcIVVLheGZR9Bc9WDpq9Nm
E3yNklPcIYEpfPshNXN6zdW3Z6761O+yG9iiv5nurhJsLa8oGdVrkLMTYfDy7M00JzzayCPmyJlx
uVrsPKx3nuTl0o+p3X7mOkeibWynHKiIFRSGn7/Y1WLDLUcIoWSoE5F2yDIQAS5x8UJ/e09KYROc
ihIAoj1ZPABX15EUUz6ZA9WXv9eV0Y4n9NbFWiWRTCE02w/XxxPnQhZ8BWBWmXthz6Ob4CYYdwHu
voiPZ59Zm8pWfZQzQULL4tWxVz21BqkMTOQ102FV51JDBYdJh9Wti43x9jCCdpGZLMUxKdmrzBE7
FbYWGxNgQWVfI9zWC6aXu1EtTypBSCbIQAqgMJ4QSIyV9XCOhJO1T9M/kutebwU8cZ/NtfgK9twm
Etu9wi9IwdWwI/kHoUsm38gVAicgxRNhMF8u+LBzCCdVOezmvPSaMtd+M0zjRtMgPpZW6piHCeF6
TSkyL0TbzIa4l2hZsjQiTuLbwsPwLQn54DbpYYiciiI3mpJjBY+0F2pLDjr4t0olaALCmOPaD6tc
/E6c8Iz8CHpBKImyo1OX+UbSvX4e5s7lrgJ5RGAi8FCg4WDsuTAfdB5hePAPnozv8sNwS12zhiHq
/dpwIu+JBWk2tKFxEOVPklEeoUWR7G3KPAxxsk4MXW4iPozS+FUv+IhjWMO9c8EMIDtyMMKNw5Ws
74dXJuBce4ahm9DGVjOCWD76aMd1yF8vqncIFL4NdtI7XO/iIIcCJSrYtZB9CB6Yaf7dath7bHYP
+tOqzmW4O6cElbz+911R0seYESsIsxDfzu2V4UiJmO/XTLjzJ29p2/b8Te91amK7EyokEeR72Yaw
iSd6uSEV54lr6DXv+5OFIQcxG3ss4kLImwJiibZ4ftk9ui/X8YZaW3JuniGnZEIX+cQQJVWr37kw
+p0x6ODmj67LoRd3bBLgnc2eruU94MXmCsRtyWkDfsu/YRc4MUXwM4KMMsaDaF/Gn3nQyXH0I6Ly
nXOsC2KqWsygrftexrjEE+tm17dB5QbpL3Z2gRDOL0bsHZlWmTK60A5nynlme8lKQz8HmXU5InOP
gGwPyKIEJXLr59EJYnAwlPggtOkCCT/7GUkLFoS0RQ2aSEw1UnweDO2Q5S+J98jlMLhEQXM51oRj
yDiCFRxj78MfMLl9SwoshzOe99U69CVF5pnNnWawxT44PFVVMSZLUSCsEwkeK8/ZyuR3DAhEBuhG
UnrBVkmuPxDYBxTJKEN8tTzSFjUkKi0cnxW+0L/7BbV/84X7elFQyuM/1spHA0fSyBo+lHR4qfRE
EXm7Wyvkbk3G9U/k8+pavf/UISrGAQDAbmbs+Uly6gZR2B3LYVD61khUN/kKFyDHqQpLKR1PIwIm
FMZgYMCYRqRYtmc+BkGVRvOjIbxMTIsDSi4EPvhk5Yhyfc3sL+mJsSv/TT+Gy+FgMVvy6lFuQagz
flr1jGXyJ1U3EdmhiOnK3/VeooVxWk/q+vDOcDctbxGA+l6OE3WnyxhcsyDobVwH7PQtojkQmsAa
o8SGIkW0xDaqeM7EGM80MgesICwfj32Bn3+Dq1yzzGHONKYL3FDtcdFtYNrh7kBca4Hm/IToj2ga
iHDlBtbp39UE1eahx5C1Jx01zh6OpIj0HRXAfWj0q+R2zYQf8nblKyTaEWH1OwBP94j1vKCguuI1
cAyD1ee3fEhyOjXyBhfWh+U00Trauk5JBuC+9G01Tnv7vFLAqnBciGES1kpII8fTQd956ulXjEU1
Z+tAVl/5ssJk0BiOymCdB6FMLNtN+lcFy03pP4p8aulTrM45BNbeKtTfY7vz39eqNcPFsKv0JObG
ZO6YSbxUvDILog/odmzFM6w0j5QDSS44MU9WjcBRUVlhYdu5f6N8Hsjb1YoA2zcMZJBLo9yNt2Ef
heWpa52ijLMF/8anYdJC1vpBRrf5XtzikXS06tfvN2/17jAsdvnpTySHVAr3q2mB5GvgHGwSy7aK
Qb9X1rxuXSHQ1/d0nJzeMSr1M8BRMPaAdza+7QYK3wph3UQFi++IpNKDz0DtOXDBbEvbGCzXJFXS
kpDp1xr90IPqZhN+FP29nNsVX3rTA7LspJdEU5wMY0imG1dHFVWV6+09RL7uFE5i7AbVHVLND0N7
xv0NPBmfnBmGVsRtzS7ZVLNjvsT0bjfdVys9v2Tn+0FMrYMjBRkRiTRP2+rHIdPrCt2fSbLEl1x+
SDC1lx6uZT/CW/BKOKcnlAIA326hlpoTQfZEIi1LfsefYAUvKZNYS6tBGvZt6ikHVDsNUZeHpUgP
5fso2FAHf3B/3hj3B2m6azUxVhnZ11PC5Ki/lvUiVDTlXxVd2xLs0hrt5IlV1wWtteN0M6w+J0Xl
Rag6Tk8exAEN9ZugsuqoACXl7qefDJqsLuHJI+8F5WnfCxplgqtDkEKjV84C1AhYwh3ebI6qIxgP
ZDpeUm3zOfu+82iceiiFbVGcNfhwJgjDMieOZNwvx99ApMOLmNM48Syc1ykEagkJh7mcmM8mJejx
+wmHraMCKqXsv6/kNxTpcC8Py91uXGmJGnXirauryuOsIz0knc6L/l9TKqv2+6aw0QTHVq9OJay3
umSjdtZuKpx0gFRQ+MvfDbhkYQAJsZOT3HsBoGWOgXVb2mz/1/vfJvQ65GR6PcG2UANFFUThbcvL
tlHXA3JO8dGlYLDF4pRGBGVlBn4wab/e6yRde9hun/e+2icfSK1L4//eiHwZNiA7ZJNO4WoiP/r1
84TmfbIfl0SlXMKFMohkwRjE5Fhc8vhfMlLOEANF0wi8NnuoLPyuPuE8q/2LJv+Z/ge6jijFBZP7
L4JHrDWKVgQYiMmaSI9S2j2gOTeca1ATFhqDZgxp5C5j2ieigZ83ySS/uJIp6W3CDS3gLcEGgl2Y
8eKFTBMDqzLSbaXYcnjpsRTp0/dkzHJtbFMMxSPTIfBGt0RdV/XIv2hHuxbTnxeOfF6qXWJs75Ky
TLhQpbrWF7ANrSioz0rqhk8qeUJriFM7AyJQKX8V4RclsRtl9eleqjjyXFM8BOZaw6U+DmT3OO2+
W3DScwSo++7R+IGSD0cHlkDBtuQCI6fZCKU8DRVbsfOT8uPFTdB0IMIRGPHr4XBCSI85G4u6AqDd
axhS97W02vRm4COhzJlHaXDo2I+lytc+Oj5Ftu6dB4c7G0q06CeCI11Jf1/gEkWNr3gM0Afw4Jqr
pkfWrrdSYD52GxRddJQYXC3CVXWz6dKJbwZCR63YDG7r0NztqxS5BhrDSSMPccA8698qBarHURCI
yCkd0UQehp6GocIT8u0Zl9uLXqSQtC1+P1AmiAD2BjBXbNZvSfOO5fDlAhPfgiKqSn6cWRX3G9hv
Ots4EDGu6irLnnAkJoRrLQYTtU6B0uDUcLvSI/1Bamlv+h5znGb85ur2ToZrlQJTpBbiyCFlZcI3
LAHdY6wRu6uIiHawsZS1f5ij2b/zqKpZQJQHO4OB8eW1MRiVmTrpvPrkPW8S5B4tWtS+jdFtRWWK
i7BJs2OZzWSsFc2ljmWedmWzSbCQ+8bmPQIgu1XvgjzB5m/bHIvFwPyIiOLne9QzrCr5hHzUYWh1
0ev0kl2jz4eYCpcum0BeN4UPB45uD0D/Yf6VSvSwZYLXFkW1C7pxHQb2hFhNLcMifD5eUV6I/rEY
qZJd2nUrdYLS8Q/UwaP2VtpagnWejMd3G9IjWc0u/W+la7vOAD9HH3m99OITIqtlOc00Xs3Te86M
1AyryZTrQ2RtfryEdHlXR+NaEyHKZtVJUIm9wH8aYbwJvllWYUts+kKX3dOyTaZrF9Uw9tvAsP67
o/YQyCRTwgvcZICwICG/xq6LkYgqY5HOpq/VVqAkFHFyfGjRvHOde8ZfKc6Vhp4Zv4B1oo4Nzg+I
XfeoBMtNlieHhpuuMmIldaycWFzzTE4jadhSW22KHb0uSeEkk+K4YxIl6tV+Ls6z6qcGxKv0hJZV
4haaCQZvlc5MwWVwDXmOPuqq0XI5xQ1k5URvrSLE3ZYPUe7fORxDT4EXpeUMb9ph/M0zhVOIvBbc
qRIppkUwu7vCvufEoKVNQ7RhH/5uEs4Kd7taNVYjX7J8dCJbPOpVSQP7Vc0HJn9q/oYxR89ovlrb
Hc/tVEdttJsf7ho5H1OJFbW53lqtXX5h0LkWhMPecqzQbCdDtyZFruKK4Ulmzz6Pq2UJqQPBMuow
/r/CyM6LV0GUD3g72TmRyupATPjkC6+nHdFlb28uqBNRJDyHAb/GQb0dhhKK4LRFRIu02MheYaSu
9sykMolVNFI6oWwrw4UwEapgXIpmE8NQhjzKRJ3HrgnwI4F9UCndDAPMFgzjqE5sMXgZB0xIf+Qd
TBsx0un4GKUX+8GljMPfBjAAWCPk/tifj1K6qZG6pFiILtGjm0NJRaraaZq4ywZPHpi55EHGye1m
PgXJpm/SGB/5wvcqYvOd7eO63OhoM0bmFqCWgBYQd+86lfCH+AY6T4hzvnexF146+davNnSicy9q
naPEb12n/cbSOXhLHnjNq3siXK4UESb1PWWxN8X5PfIGU6aiGHpQ5YHXozemgFGbhlfVV61DtqBm
8+hohXX3SHAcgyHsziAc+oTtVL5yaqnqWQcJX64yS7LL6jOmoJdIHTef+i4UWqcQWdfYSiA2rSIE
U6q/ohD0NDFq3DdFRPq18nQzFEzAROaboEXDabpt6R+G16Aj96LAHvjYPo0SfnP9QH2kRMOBJ4IZ
vreREXVfJlK2ekXi+JUbveEnfSkG9fKsFDRWw1JLIlTxpnlfR3v4jsZIWakOWHNXsVFQc4sun1Wg
vYb3fe/iIDhck4VtYO7Lz4srP4snhTXurDh6PhKxzKUzBJyGtElerGUrYITtneXTOT/PEkNcexkk
QZQV5ub9qCGTZTYKL0IXZUlBvGVZJHDGSAl/cd3CK1YuuUF9SuL8UXVPIDtZIKPG8g/ZN8dAZLwO
Zj6bc7u9TopplSqIFRXMazAFISn1EHf8xk/jmIJeQ0Od+Xb22W+l0agBgKf5Thad1eAKVWGYZgXZ
xiVCjjC9LjQFG1W7QFROYyrKOOEGKhfbIS5+b/8cdnoDYXqr5xgdonobzRvivlLLVR0kyhYe0i8i
YT4QJKogLFLoy5oGzLh7RTyWV6xvPKNNEPfmiPKhI/oxhWkqgl/srHhG0kyq9OTfzWEcz2ifG6SM
8Iiy5eVyADq+moHuwIEuuOqP8qOAZapK8wYoycthbbXGlDgxBrieLlpPFGaAxYKY4F2C6aVBiD0n
eG0cuIN9S9RtGfsg29TR9jZAVfP7iwsFqm6sCC72IbCr2bNXLfH5rHFcVlTgVqtvEe8BxbcMYfIz
FTj21N4mTNNtE5MZBTynd23aPeflHwYoy0KdmIVqDhrViumvQLk07TdF8+LU/I627MARdEjZA2ZE
LIm3eW+DSqglpb1Ni2EHMEZVnvQIfTRWQgCAVUesw2+M6bNesIzai+sCnrNZ7/tBXfTjiMA2coRo
ewCkABo6XvKbcc1jzV6yX3DxArvmCV50F4eBmdtcOofe0wE8bxs53efoZ2WC9x61Lvxbqu+0dLRA
3tD8ctSIF2/LKNwfdiH4doIr+pE4UasZQtW6knvStDPpVKKMVg1vYFmZgB1eFjIOGKUWCw/2RBKn
QJALCAMeBJ7BrkZYMFl+qR0UvOSABfyTnqJffKfZ/k2DMKwWvMecXymVN0O9PvwhEJInjG4YX82Y
nTYUHEE6MLUeuCnmFH3qjtlzc8NBRzA+g9UspAdKq5CPO6aRYZbC7at68FJKvPQo9vnBhr9aOnI+
y0dpZhh74eFC8Za9TN9kGqcgzGvHwErgXD3sglbsnSfbL2htTqjPzW7Gt6alFf3mmzyZjoy6DX70
UrVxiE64WnkfoSPqEXSSplRwQznJm9QvgnM8Bpn7g+GZvALhSMKJQpcIeMMIYMN/Hf3Qt+pYuhwj
LYSB6lqCxWWgx//+vo+pw+ZfCW+j1ZEOXQmRvboH5D5n7A5FjbTuGe3sLu8DRG7BeUNlJ4UTzofV
DSqHrv2M1+FKDOf83UeM1iHJNH/tIsHQoijoph+dVbH2SqGCEDwFqtBNg19DtDrdz9pXvXYzB/JI
dZxX17IFCw/7aEfT1DKn4/luiaKeu4gXxsRElZaz9aEFAmcGtHUwZ/+fBfY1Opibx71Ad7+Fjlwh
CDCO17K+PAtF62rcyLtNXQta78ILLrDFRY4UKFjn+oNtfHkUIVJBtQNzV7Z1ISEUWJig9uzILqxX
WIIaPLCLTW4GSE0VEsJYPLZzJoqSpE3iVi+r1jvp6cE8x7F4X0ojr7YD9gG1KcoXh/ClBLfuvOhY
pigODOFnqOzet6hBpZkJqb1WO+PRUkzRVYcbRRd8V0qEK93H7Oe4W2AFImCSJ48OYmBufVjLYq6q
HAA0jfX7vwKxBDgIs03DcUN1EgYcauIY2NA2c/pmPBUpLSmoDsHfZWmuAZaMww28BYv+OL4xQwe0
VTjl+VbigPpTVdVs4FgmRHOZ2WoiBdRMfyJQ/mFmbLc1aIkWi3Z7lvA6UZmD/UUd1yQw5Fr+oXDE
AzKYnsufV384BLeXKqaH2lqmnSEk/KA9+f2HYLkmQybDY6nbwUCP3G0nrWGM82ZHbVf7zWscM4wb
2KLUm/Rjiee0eCjW0Uv8HRvFEpY/JeBGcbY0vOauETj7E/S+UZ3ia7K1PjCk3Bnk48hXCWKONHDf
vLYHG7qGvU80Rrm+7y1QFbgjRQbiJS1+qRDZ2D6zdeR11G889gnoF1/bWbzH3y0UqP4ilkMf34oB
XB54+icnsZGYdvUYf29Y4v2lKzaIuM4E3eYq4HG+5/YlbJCPfsEaI/ksNrj2jZ7tkW/h8LEreW5t
UqfukA5nJpkh0HCQUmKJP+spy/sAtFkGD/0+pOPcxPLz2Npp0Hf8CRCncgrpSA8H3xsq4e0dPYlW
PJj9wI+wRrk/N2hClCctQnVzPUG0qCmWenORPZQZ6MKjCefwn2LbpBtb0m8zu+sDSMlvWWv+lxAG
tojaynDUiZjbwEH2wOUdO6/f7MUkJX5lxZJM5tLxXucw9j5rcXBjS2KktQORNeq3v5sjjLnXLUbr
TKKzbSIWwJzrh52UGzAA00zwO9s4A4XT+dG3WvuP31UPYMj45WamrzOJr/JWs4mrxhCfqFkJFvxb
97qACz66VAcLqFvdOCq1AKM6XEYw3M4jLyN9JsAYLwFk/CDF/nrqU7KRcGk1Rko5KmGdEyaAMI7T
pstd5OZlIebMz0lomrFz+Exvq0a2xiY1xqIbGUNv+WAsFlnkqNhStH5e7Nv8W/prIBiS2qqgmb9C
yTxh9tZ29nq5Qa/WiPCBxAWs1PEojJizBJuORzfkrB728qWg9ZjpbdO1GidhxrbHKyl2Qd5TalnV
H6tVOcOBRcuz5MuaoqRgVnvZmK97ONT6qYrIkZyNrsfiZRJBLystzR4+YY7AegNCKjAcmGv9kIgZ
SPhU0dUEctSMnTCLD44uU4vPy41cR6W8Jgyqf9OtzysmJe6Ck6Aum453qttWVebFI2wNXWaZMC/1
o8HE3ArIifUq8EugyWfW6ctD6VrkLfP30K36XVTfTtlajrQmdQ3rq+DKKnd+crif6QWCW23ALK9r
RFEkLlC7oUQDgerEw6Pidi70eMEJQcHBwDgH7vgsRXkslqxhBghL0RkbxwSlV0TlqOz3Kq0wYyWR
DIzQhRCrz9ImjrCVOpv2NTbnRkbkwHpOl+/jTPuHPGo+tn0no1tH/tkVahf2tlmB1Xq7Ix4wrdh+
UJULRvMgz63rbDbMOIfwBN1SITuH8m7vvVmEjbRUucGeYi27ohWmfIKuaW52sDD4olTi7mUwIQ05
HzVgNIdLv2lzZk+OPfmlL96SXdWXBnvGGjlv8g84UC3WGse7pCJteuyb7el3ndgn09YTatEVLlVp
KtYsQt0KZQEyTCQjHuye1mxB7/3VRltS6nsQ7ZSupkS84gKUFXpbFaABnwz1KLKmNkpwVTnLMgF9
Ika8kOwMAT+ApwOXqy7qXtmggetIM0p1uMmtGT8O1A1ES7FiPS2SOLzECV8iJKIqCwrFXFebW3Bp
8Xm8mqdhpeZr4kmpI4/jtGPlBdXk+AkIfEzlYEclX55cEwEbMxbes8xJJUFz1bvg4zVTiotoTiW/
xoGe9qHChFLDwHXfk7siwwGMwWTpMmErwAInFWEZ4vbMwzgeET15Fv7h1hNd+HS+0qXc5lKXvuG1
/IoDKoX1wbNjVkKat64tGUpXIz2vtPrEvTqYgiyeaHI5GSb25q7fEdPXCbXEfR1GewOb1Wm1S0al
7xQc57ILVCmKavhHbGiNXDnJ8WMj7VNv/our2FPHemZkRhTdGv+ykDBC1/OyKGucyTeCcSzu2Bfg
AoO+E3yYE3ebaNgNNqDhpANPJZqjYptqyMXDumgFgjynJMfOi5sZsBkNEatc6Z8fwcm3XKMji5A6
oVay76CWTLZ1lh4Yc700N1UQT6rp3+f+8c62cZ+WXFEM7KLWJoADiDplGaLAi5QNqI/DpMu7+mjy
Bklj8ic/yp0zK52L/qMPbndRuihmVJU+IRtPRUgxBAaUJKuOsCcAZMPR+JpwHeq7cFunHh8ZHUTq
+Hh78BikJFB+q6SWJ6VY3UgSE3+VvRe8lEZsle2stGLS77zx0tnP2AKW5RFnt2KnqfFg1f9AlAwQ
HMEbr0GJOM932z6jsefssn+GSGwDovLyDNUoOQmqFv7gGeGqA3NeS6m2qupxkNJicXRjUkd+8E/y
TPMJmMlusbqAQdR+0jib795nAV9bugMnirtJjMRbtENOsSDYsxTVjByVNvbPbvgca3DDxftTIEe8
Fsw+rmACMFaW7K2DDHi6XdwOeqgi7ADD1WTqPceXAzJ3gDkfLF3O4fUyjDfhTiEV5I9FwkQ4qvJO
Jnw4bP4wgtQ7be3LB+6C1QW3S16jfUU+zMZUwPivpDcIWvXhSLd54pZ3PGKdJuyrq+oFjkKyK+rI
hnQih/5ROww8jxL7q3fGWwX4D1gwIBSwvyT6KywBjf+a4t5JjN50p9D7chFiyTN6L2VZPKkWNaX5
IMPyRPab2Il4QID3JY1DNKGnEeVe/5bFfvP9KpxePnX+WotgjEYzrnMqN95rmIXCcCEMnJNzgTxZ
6Ad3CRIaoiCTT7rJ8W7MsqK1nq+GBs7xgDo9MDUfjlcpQvLbCddnhihO6e9BQZRO2zbXv0EK2f2q
mKdgHdRTwfND3JCQ1Le2fuUAfSN79bozxdYbO92dlBG5hjXiSr/jP4q3yvl+4oM2z7k7yqZdS4CY
QCd7HsSPeJXDoS5cq+Q2g9QT32JjrEUIXFpU7C72nJo3ioLmZgXFv3xjzgDW0CHSsJWiawgO9oHv
sZxj5JCw4w8Us/4blx8uR9Cm01+HslijA+zPfeNyam5Pk90mqoev+ZYnb6GJ3kpWb+ayYFQ1+CcI
nARem1b6sln2V7rtb5SFdMCxKUJv8w+llwTNwtXjwnTln+sbXJvY97k9qnLOHCXZeoERlnII3fqz
3SZ3T0XZ/diQBhIPZvNyW3wHOnqItWHnu/4Kv9oGd2OAGeQm0yJQdhtzFY86zLvAEpmYCOO0cUeY
Lj7KKeFQ+SmQtsJIc0bICF2isRgC5H/3YdsWq0rTubnv1cZhgcPM6+Z2lIlPI7isFePNkIxX6bn+
J2N2RkAs5V+9GjY+sYlV/0lwkhsrn2wRmWFlpLGxhVW8lEDVdLoqIOmnYQ+YICuzH2p9Xn2dVm0K
Dd7wyBUfJ1T9sp/xaLfd7MLenDbQhzDWQDh8vAWB2tH+FASdjGPhjsgvLQP53/cURAlxiXZtU8lN
iRbs0PUlMAKXItuTrs9D8bKQ61mtEjHndkMpFj14DGeBpkhAcwb7nHMgbMSQjDujtRjB8OAlCdG4
Vou2G29jAxN8eFOC3gp+pFbvASeDcAwNZgVDNzBjRntlqqmWFeVU6rUlCsUOUzHo5qh0P7mZQbA/
7cnspskNjbF5ecAFK44cY6nMl0J36vsodj661iYdOCwyWgzw9poTugvZh+fe/7SHvmVtfMZ5Hi8p
kBVjmW9r/u9UlXjYyxMSEVLzXGjyqMAZihJ9/VEr7GWy5qYe+oVlDgM91MEQQupCRa22yEH2twoW
wKq2FmkhfX+PgsCD5qw8qasyhIqHelHqZbcb+yJ+bDZrufymsZXrqovt9cD8o9dODRO4vipgNxxy
PaGfsSuEGjEA/ebpY2ewaKOor/PRvMQDPRwbstyjHOsq+Cd03Fk2KBSc5Ts+SEZife+H3gWACLp9
V2c7rd+2Suf33mSV7aUlJK0P7Qqqc5BUOi3/83OhebJpBS/1b0mim017QxSCbeZdqPVxyQudf/A0
fPqGcJo1+cFpYbUvduSLl5nWA5zUTgvopikqlLZeFYCISNgfebtTYSlDVSTdhKFNWQm+8PkBZ99P
OkRgC3ywzLptyNHb/lLM9ZHVXth90B5cbJ3P6Hm2flr2t/Ha2lvcD2kIsB1PAViUe1Vy3wR6SZG0
UmliYm679zQI/7UHoSHZgG5s2j23kxZ9lxpUh3vtLJ5HwU/fxNpbtXYS1eLflFQ7HaFPG3qHVX8t
dBVGagVPoVlrEHPqKgfna97tqwizpayaiH28HnczOWnouvQOoIE0ZXxS8sHqinYSkNQjIY97e//M
XRk4bj4Bz1E/n1qbakpGqSy9zKNgYvW0JoEL9AHB+jmD2sSLcUetd7Gl7XSjteHvmgx6kUObidGs
bvB5nWb5Jh9cxX8guzkHQxiyuOiiXwKTBaeiy6zzlatiyfZgo3b4OUGJspM14sMjpGF7v3gTGI+K
jIV1MJNwdZcHHgDwT8AlclkUFdaV+0uGqTxWSYkCcgXo8xGeTpH7qf9jhrKWSTy3skrwtANysd0p
gSZe81jDoYKZ3MGyzs2al3lPCYfE/bsqSk4AhmX4H5phK/AzFV8pm5RM4k4QZ8QWZyd+QNzkGnSx
igUsi7yKaGKszks/RaAuJ7oGSVNcQzuxcTl7nWqmWAMcRPpk2qTuatdqY+cBUdDdUcUeksUHAhLK
WGem3/GZi0nVNtWfQqJC+29swBkl8sP3FDJnYIkI1wV76u+kC69rkTRFSI41RdoGnSbrkxCQ/Agq
otZFTt8gGHVtPKHUXBqfPkSblQ59ACliv35BOlYEb86pzjZpBoZUmGSxW9LbpzxZAZJNLmEdUQtC
LYF5P1uZxpVDS9Uxj5PFdD0/v20/Gva6WkSA94moopgAGAql6LXtH1ppzPXGdFcXbKiefNY1+Xsj
OfYPFX5d4y98RLGVAYECPXrF3pEX39U8ZfyPGfhVoTlD2nEnVl3IHvlaNKVaKZx+SY0o5Y628wUb
sS8Z/K/j7q2Z8tWm064PAqw/ib80/D2+tgwYdSv/FueVlo378RyTYHPshxSuwbSocwY6TOBzbIyB
SbWNuZu1BNxHrjedRo5JhD3hvwxId6BrfcorpZA17B/AYAgkiXKKHGo/guVbhmoHAjt0Xr7FgReW
56Xv2LAEI91+mxQqa/ILNaN/yiWONObnIpd77ZOaooVQy5J0sYug5gL2x6lzkY2uQiWVoN0Xy0By
jobrSRLTdc+UOA0OlsNxzZydp14zkchCXypqLZ9uP3aW/im1ceihoZj2dc7Sw6eClbL+KVRAIVtk
rljC+hkJars26kdn41ibidC1+ZtPOapDRyGPp+W0akuDJzhYS5CI7qMLYwRI62xkfbhSlLxEfLBO
3aWaN2GgtdXWh1rtC22ODIAsSIUkAIt1IncWwGqi4VxvA/sLHjB9CA3kIrOYgw5yJXJukX20B1sm
YqdglyQ1Q9XEH1wdORrwpSkcSSMQPeWXJ2Jnf2yOiFSj0GyPWNu+B/9mOtcca3cqKoyTUKe0P4C6
jnQMEXjHX09tvuM4h0CSCaisA1+iEvFjFWzAE0Dl/S9vMtZs71+4uZRxKRuG/JfCHyVqLHwZ2LZp
200SNmsYmPN7W1ljlW7Qwp5t7a4YlJdOpA5LvQsEyo34aEXv7ajXG9qCcEddQV0dK/pSqmlHWNUA
9fTRUGCdeDErDLRiHqQp/MO3xvPaQuuP4Bl7F6kFNdyLY+lVOPWKpD9SH1ptbMPcL8zUaryxhlho
VdiRaC79SYu7/iF9XSPrjzED9oXbiTi3jNsDShHUTYswVsI+fNPJ5uunZZaIL0NbvIUt+lE3WUkQ
v4svs1avR7pKdtU6aw0pQk7Wrdm7QWFfQGqBrN6+OVsHNn2yZ8bVz6DjX2cEEdBph7cgpt0umcBi
FlgWHxsv5mgJo4YOjOHxOWi+rffcvrUtjDGu66UhEig4H3YjkJfd1lStB5/M2afNVV8JnjIOTBN9
FjGe6rlEZLcr7p7/WuLp08zB9UH29PpqbfsGUyFkl1k2DduaSqsQPqCCod4F4PRnTfweGtP0bTej
GCnm0vtA2DOCGNFi2h/irHQrT4+zh1KIsUPFRwakaoPs7hvXCz+qQKWps8+SFsxgBGcg14Q+97/v
hBdGNga6KQoJQnP8MAZIzxLAdIy/IUBUo6XaL3gt+9t4yJsZvo5GqcAIfBUrGyFCw3Ia0NKNcfUo
159/sBfDsCCOFDIhz+pLQid5lPUdxuZvS4X23DQN800THNuIqLinX5+9vyp4Rird9clvEggZeiEE
81tYnyiYhmW2Z5zL74nuqvvzhT05VrgQyYzXcs9DEcKmKF4QKI/NvxYLSQiHuwtksSRQD+AjeJFp
LC26u7d/zHUkoHK7ZPapHAe4wWbuhXL+kIDphryhN9bikuu3Rf3PJ4eUvYh94iMpYgFm7DyjHn9+
+OIz9R00QAIv9UfULtbL4AFYVzb65sq5MgZNFXOdhB2eWHRuaelpIlG0M5f3UF4CPx/gWBq4FfHP
ingVwDHxhABLarFGFe+vc4JW4wBoubNCizm/U0XRg4SzbmzCInJxqXV2aifEY9TKaebVlfKqNbth
CW255vOl5TRmqGmVvSj01SqD4DmxTLIiid/FDEW02cwhNB6TWxwtSQp3eRpU47HIX5UowyMMtJB5
1TTBlvkvWphTChtYfvS72VSeMafVfHs1uL+Q0GN2JJ9fSbwazSgrx7ye4VjOOUdW4Gr8D9+pFmSq
tRkVDoDuseJf4z0I6Ik0EtZlJ4kONvLcCxUGvHGA/F54f1Eo1AG5MqR7UvsZBF3rHlBQQqFSFSdy
XGTMCgmAV7myKOWch1nZTgkObgeIiAiX8AoxZOkci2lkqQSt16n9qXY6p4wjxZPu0seCTb4UuegV
lhTmPW9oDQFvcOM1yQo34Q+Vip/cbU+aoMOG8dtoDjhdeg1UqrJXZiM1J0bZZbsYqQSKycqeokvM
sVgUygQSONTDRpqqvpC1NcTzYvPoHBqBT1sqIMreweYw19qpa2ScvXYliyjkei+OelMwKhI1gVi3
XtNM+ww37HextAglVrJwshtrds7L6BFVn163quQQsqFuwKIVd411YWIzHUoazToAsh8aLl0OKDFG
EMPzXUtzXeglSBpy2xRikaVYlTJeCF8u4Eod4VZDzE0DbAPxzv8HH/5IbJ3jErW4R+GsRqZNvkjS
0nz8QtRVBocX7kJ6Yxm5A8OBEBjZ5Ux3zr5nEpFgWwT21Mgh2siZUaZuj9Ddv8B6Cs0D6SyolciL
r8aeQVW4pzmxYmvcLwf+xJBgeMcCh+gtmU/UbM/9glnenpN/bqZrXNLiff2+HohGfizeQ/ixkyup
9UTle39OY+DD3Xmuy+LHR4gQg8s4lnY/uV04MuBCLywX0+z+QnRjzrh1pyN8ujEjcMQjhaOq+0h3
GEtMok5GeIdxvZBIqgGuMSX43L0WItRM95JWFNCnv/KqsML4KT7gD0eqbEdPP2+2slYbbvRQzd7+
7QYZ0j/E+Qn/Ejh6wLKfw2lhS29M85fn0zo1Mo3ntEXxX3cGpvt0H54KnXsQ3LI/72vTLvToVEPx
Yqw+qN1Be3KS/OEuf53A2a3cfUC0Y2bNNJoycSL1c5wBWnmF74IRaxa3DGXL1ccDdC2jZ18vkboY
3Uo4a1WG56xPV3FuXLoLe8hODLgSKJt0RA70WSMWEVmJKZl1uYUyYTOpsvvtIk5VYj4/bGKLnL0D
uVAZvYxfZncFAkJY+cK+1McRmh922eJlmXJF0q2NhYKkKvxSxZxHRJqbo6ThM5Scy4qNBNPoTE8U
doRxMaY3lBC7+vKV9fhKtbd9TcSNpHgeHyK9L2TgPKGRx6UTbnFqUgj8rAtvTMokdaGqvxJOua9w
HeAWQVrtsQEpsRdJrVcxdtROMuBUen6bn1e0ABzRSLTRx2l5UStOH/sQKYMn1yihUVuP21zKRE84
qzy7dC7lfKiVtzCyfPNOdAUQDXvneHVOAU/Xc7Y3pmAy1NFMOQ6dtG14q9BMSyKA6VKVUBzxSEch
uARKvZ9LssVoXDu9soLmuSl8lB7jnkLUWLN8J47zra+TBOrQ7ItZP0WSSG/GWiUgHKARdciPuU0p
I83pCDMB6frVRqpZYYGrO7DyLq3WOCJk0P5sypO/o1Nmc2VJD05hp/dNZJlD3uUHGl9uc57zgh3R
FJWHyZD0Kabw72PuepN6u5TwNA+UHw5A+YgOGj3WoCjd6t0g4RPzE/lLgOnMnT3oRIPmIdyjMLC/
Zw0eccD2OmqSXMvOKcpsE7zb9lU96qDd5XUwVclUjKyvxVEviXn4FwYroF3RFLAzViKaplxpvqti
TSgKPIxK/m/EeD/DVlVCEag6LrV//DNzgH3WnlHXZu/1fqUjU2bHsKJu/IdMLtmc5HvWbjcOO+KW
wTvKCSD2YNxBNDT6lowSrNHkMj5yfI8SGRjJlvBbdji8QFM2RO6kAgo3MFNndHnpmhCjrXMwIWf6
2PGH4eqUVo4V+9vQvex49NEjq+AfxBSA9+jURfYlB7YMg1Rmb47winA61MzaoPmbpqIJraqjmfey
wqtIwACNJd+gHuGtH2XUngV30Sg/uRXpnxWRjaL+5aCFdjH7W9E472JIBSLzLxYumM9yv9qrmWQz
qEc9P3SHmQeJkbb6ecMRci0Dg89l/BPsuXUon/13EDboVPxWyCmOlnXot2rHkPCiQEnzCNoO5sCX
QsuLOAUR8zs5wG50I996weD3l0vRZ1ieTWCgLOiAc9+IxK6Etobywz19tfUZKx68o1j7601qDR7n
BnCaY3l5WdgxhJHKaspI4QeqWGW3dT3Hga8GXsWP/5VcPOWd8fkqVHWk6aB7EkHGviwitPmoM0Ho
0sYz20m93GRHxFA0MeKpGNrNqAVlQAJJYjg7DcpK9IKb1RfTGDCsM7cYEyarXOXWoqZbzzfYa54X
fgAChgShSMtjXLsRaqWgyLedfOKf9/Dfg7yymRzaHmQYgXmQya1Kbd1KtnI9xZhVuNFRc2tnu6a0
PorBK+N7Vv7al0fTCueo6DQYpD09EkvtsqcbjMjlAxAz28m/e4Clm5QmflE64U+DfK6f8SFn2VOP
kxGrIOQDcp4LFTXqRtB8zruWMZup/LGNFHPoTtuv+wUEbDe+9HnC2x9EzvYe8pj2JihK/+5l2Q4f
5ZBJcufpDJ6uVxPgsrzY0eiUZgHkSztCs0Q5sEC1CRamjTZeagZaWP0CRHOUu2m49HhQXoXc30+2
ODySw/T7pWu9bmdhNWi8Z3kl/OykNxdi/M01UyL9bSTi01VZtFD70y4MOUag2pStKgkNk5tmg/D2
wwHmXaf1KkqhPTSv72ztBY0jaJ6kxtI8qCw9wpY46cT6BG/lkwqZpfhgGIk2dqGKPQcT+A+lUHHg
T0NREGEWz4ZmAmKJjnHfkA3rodPpqmTB5UsvwOydVpqsP8CvX56WDHySPQ94Jc9Zo4Xl1hb7lBsV
LPXrrk7r7aQwlpTCnUlSa/1KUuOLBfiClLQSMK9ZAX6p3C7ZynMrJX3tOv379OZd9Rn6kBmgWBQy
MtrFTEkLDuswHg26oEFyiy4Djo04VqSJaha6qXlD9VH7btHU4zpWQyTokk2PU5lZk2kHVEL4LDk6
NQkBLTh6fwMn+Qr6QKu1BULtEyn+yqghmJZpgcbq4JFnM0fkIQNdy81895BBgPRbAOCiAT2/wPpd
A5Ms/SrWNTx0+4JWi2jul9TSR8SvNffgMuHIYIYpA07EtI6j93qxzP1dHCLAlB9/ZZtwz9pus0cR
hRq8/FDvpRWYPEDKlGPzV1vatLA1Ksja8BgP1EhfstvJz7Rh4mpCTJu4zQ78ZqyuUNNmaFfhQnN4
FKDQU4awAiUeDYnkHFrLyxkFIWSe4LbvB9rbcbaER0H2jicuVVWdIAyP/oUtYWs79nE47cHH8iLp
BqpXTijoawwbM5sn8WmNLdjUme51R4WkJk++TelGMtyb1sN8fIekGHZIw3wXtLBR8p9AGaru6xwm
La0xqKrrEkAX7/vLNRvrrbjyIdWLcz1xvdTlfUP3ZudGefhgEYA/RcfTLmZ1FSPPSgRIuAOIM0XU
7RkvLd1FvJxQRB1NpnIPpKUzDM6ASJZS5RYtCVkUy4QQmI0eTz7/X1U+xS1T75cQ5Fo/DZ3x34Ky
3p34cPhp7qHetAreIP99JVKt8hRxW9mt4NevwTgwb2ZhoGgSIMKf1AJd/UaC/AEzqiQ9QsSg8RPS
ExRcMcYVt/wAkuY0totbmIugdie5pa2Z8Dpnw+MarXLewkhG89m8dLNyDjQN2ny2QKBAX3vPn7HS
VYXtnpS5YzXeDdcQYUR9AzohxeVF6/q0Mt8ypEFyboGwA3xTtS/0Zjna9NhFBz4a/oH3mIa6vRle
2LW8dJfFllbfl1L88H+AFMVIMYwYPMvS9Au11V9bwa9h33pRCI2Dl9p59mZqzIfhwiCC+9ENnqQa
30PCTBnezvJNdTyJqS5IZCOtgddjbCWz1lex2nu3KDXATTX3PkknzJ8seTGmVQW/qkAeoMQDgb5Q
bFObf3am4/PHZABQ4t9WsC8B3bfPEnZIu9jvCUYitOaurGfQ5XWDQg44KVKUWGt4c8jezZggn/7D
yfWmcYCsl5hW8Jr6W6wwEllQGLpd8zrPDJSqkhvlWm2QnrZs+XAfMThO30FI0Xa/rgAPSxyLBVg3
1zve/p5MLlTqTZEzg9d2tVh7Wy3Ji6ZB3TqA1RqP+avLdDa2yxfYqctMsvl9aRiaksqBmU7GI8MT
/Ic/7Xht4X0z+MN9DyQk27OxAWFLkgn0WqKvOnHcsiQeoeqDrXLKnEy4waVdzyWQIOgl9sdo5faf
+2UEiV/55tOjM1UbyLW+K6A69Rxr8YbngQEZ4i7EIGHR2zNhYvLKF9tTLLYu1nRrjlAxvTqrLwvv
sZnsAp+HuhfDcFhcw/zcxDoEUNn43YIeLKqcJrJCk5FvCvapiC77mo65nokEwYGWlCaK2VynOSlC
pxqZ0cSfwJBv3GVVbHXOlBLe33WsGiMHzzZGfyu7h7JdiVoYomc3IaIYpWUGpwM5nnGIcrGIob42
d3JHeSXfkC8KtFa1sa4fYrejDNRjoDkZm+SUEgrEKC5YLpYUxSuOLYucGxJ4SP6iHdG8v7TVEFHG
dfjsdmQpTar4OMUyfm7U/qslJuaqNbrfD9ooWO+TuTijGmT8aRaoy/XA66RwZ9sl6O1AE37TuQHa
UXeUw7GJ9d6TldK34v/h2VER7GqKulFWeCcrBZqrWSSuFik5CdjSbtNurIQT5KcQ0+cRXT3QDBQL
KQO5W0+1ojg1C9gwj3aGxhDKtlk4nwhCf9X41IQmrIEHFtkq8zmN7rPDCI7QAXacNfGGNYG6Q0/a
g79KT9p9siyX0Jzj7h14hgEUYPftwMebnIfgqUF7EnPy68dlZo9DbMFAr1BMOPeRYHCFgNX6i9Pe
jqQSkbMYybTNvdLKZk92wos6xKX50ZssQOpm1tf+lPVJpu00J6d0kqWsV1MOUccWXedGgAOS1Gl6
mEck9Zppk0jDWO8xA6SLKCCiSAMfxCrHKFFdML3/TKaU1ZgNUY/1K0lf4UGDISd4rvqmIvTQgpCA
u9hpv6/57VPz5O8Tp33jSXu9qF2vTV9YkjknJNJI5XUG9Em3Ma65Z6Zh0YV12DIoMJd1DAeC1WVr
eah/r6O1XBpRLf1VH35KwBC25mw0yWN9HCvqMmF/+lK8BoAOB0RhC3lJJUGJXVcQCY3o5MP8JvGz
dN8+ClXS3T3+2Jn/taEr1bgUO6+yBgqhXacKb+4Fr5y25uaBxRvIPzdQZd1vFAv/Ykdx+NoxTU56
T4i62f8pWK/xSMIkWwk3mhjdo5lJZwed1GWcnPw9hq7KIUFW/MUyPt018dtucipeH1uuk84cFYc5
zlu9Kfi+/Ug09knQefynrQ+qNMHG7fCiPrsc7xtc9aDKh91/2zV76RO8Anr/5h4ZGK37yaad+Cmk
aICg//8tGKqNUg4VrHk0G1qzklv/r45xRXHguhZIsQ6uRhLMh4lBdle8nSkyaGjjqnEEuEzk/4Uy
OPtjeJ5dbHPL/AtRtSZfhBod+3dmNvnxY09KFkIhyuehW1wPoDeIvhs5gBh5ck1LTP/Rb5itEeML
lpj6Yj7xv0ADazu8EIsAzyrYeJzxChF+CduGsYIF5qUsy/YNeTiW4fIeFuZ5hmnGyKnbMn4HidrE
NqnhrC4w7vXbvWXs1jXqB8SOOHSIGGpqoBC1g2TLXkDSYSihmKsW5wInbG1ErRKm+bDU/BIcaAAk
mr87YltJozYzhD+mngemngGDIFo2zAWTFw07OCfiq9GZbgrLFk/Lt7lpwRCXaoVdudhyp7sjJlNL
N0kLxBEVvwB3Z9C+eEkyt8BMCcy398egnLyX/c4kDLY1qL6FexXvdMqVjcQWwN4zui3et6QP4LJN
9jCKoHzFWGJE6kl0jYlO3uNXwy78eyzlq39HGlGwvFbEirlr94HZgWGfQqg0p3SKOKaXU+uW7Sfw
CM9q2Dimn0zEeDi7ukESfcrohSWfgYNT26pRG2+SnGe9T/ZhT1j6rbwfbd2RVI3tp17E5O2s1Wvc
rAOnR/X6j+ocOXmnLzR3nd77MwGlxGDg17B7ipJQRgntjNmYeTeUgKr+3sLHbRoailnx2KL/nPa0
y/deryyxv/xcnEcWKnn15iJUt1P57rXxeNaruW4hOG95X4W+ndyaraw3U6ioOBdjSYEcIO8CrGTM
LbuJHFCh8ljf+3RnzhaOPQYquqzbz0V1GTW0ZgM5xcfQ9BkqiP8X7y4+RjEboVn0mVieDoUUSR37
/ZCn1Km7CwYtegxgrECUmTl1vWNN8B5pIUdbNW663S93dpEYsrfKqVN5blTbrFACWscgQTmSTuwR
lYvEyi/jBjEpCjojR2hbKJM/RsyAvVelKPFUH3w2sT28EQV0W4Jw+K6j7S4QI1q99anvL4tASAsN
0kwi+dP+ibHSV7SnLvGx1aPXuZEBNR+krXApYYU5WST0QFdEUDukA+DCNhz8xjp7QGBhsyb8Z2Vx
ne6rh4+J+V6UbeEmyz6++g7MTHRf+NINjUi1L6Z38y3o79tS0HtIny6LcPPBlSjFHO2RLjQPV4h3
vuFx8PP9Cp5CBeK6q0ZXf4VMXH9cKQiE+y5+9u7wP9K1i7QrndCA5NeUYPjhgze7/p6JwDxSoYjx
vrLZTbp/LcSKCoAoEbPR1yqiwzpXz8xW1c1YyYnxv7TrHXn+KFxzTbAU9EFuJztyk9gtkztyCQyi
I0fZl9v9qE/2L2k3o+Jz5m1WfAMMPJEGxHoffOHEnIFDnMPHO8r04X3qW81TD30jUjv4cONe1DP3
Z2znQYWZHr4YXpBrsZc0poqa6bwYkUynmI8+qHz6uxUEVOOTqLitRGx2o2m6BJrj5ClzS95+kH5g
pyU8EbQkjga7Q6/xfE/mpiMFW074WzjD9YPioofPbayH+lUuY0mkTYs/ucZXcDrwmyRZiV79T38P
sgUAcLY6kaJlr048ei9YhXVN9BXVNYZ0/GBAAU5dpMkpBbBjMF17wrGWJiJvbBQ3KpfSvBREBQgR
inVKhFkL3kdUkot8tdRgtVpbZw6bnmW3GGGZZrdHpIx7+Bkn71EW+EMmFm49zsfNXY/yy4pEOK1l
NiJeXFU7w7/f59BsTifKoaOgFBgMWBHNWBL9mQP1K2qEj8rGtw9h6zlijIsgFjZ3O9wlQzUQFq7a
xQDDOBbnhbMM8zGs8/CxcnPaAA1DdMwoFD4KCYxDYvhuvLENGizt1qIQ+SvzdCNp+iH1mQOc0/2T
3FjHg3Hz6Thw3LUyGI+OR7g3i7DfTdLVetLFb32DRHKez/QMuvAGkEiQ0eVPBZymh4uCVPU2u6vg
lLf0hNrYZA9QKkv4K9ihaf+Mxby0CnICnmeNhTIpv4gtkzldU+xFVX9gl05DRtv5rVIxoByQ0DpQ
wVa0fcLwhkbbVZpbX5W7fw1OSqx3yB0TAdUl9m4EKMKBEXVPv6jNZHT6HbqqsK+CY4o/yH6FQHcs
FpMCIEDTVPpJi5rLQ69Kqp6MG33a3opQP16FPAkD7NEDN1UiTaY4oLCe3O5gGQNjht7XcxiTsUdM
l1+aP2bQyfZXsXJQ3yhUGMOhj0hcxcFw821OYuI0JFR6+bbVhQnH5hV6VWO9iufz/NPySQVJ+9oX
pBB1i9XsrBysH2HtXHSe9YYkfkJJJjzNzf/C5R7jcDq5J3Cd5Kg6MClSgLQaNX0KEXW7SNA4BNV6
NXYmpNTBixqA8PmHQhZFhkEbT+qQkthy0jBq/A0TtyozqM6UP2RAtv5W0T6gQajBV5XLV7FBo5mK
q1AjQ/TPP8JTT7u39Srca/kCHe4GuLVn3RZRSrGORi9uQElcHbbAsiC5zhYxhZX+KkCjJeY76x0z
7kU18mEYwfpgS1ckWkUZ2ey2plrDbnN8pa+2tbiUhEh21+8eEavRdtvL2z0d2q/Yo+3UDIfkoMKp
/rx+e6VEopjU/xVoNLEidLovne4g8kRKtSB5ijZ8rIa3qLZmsOs0b+qYov9o52Nw7TyHo6ENByDK
6CD/+sXWVngnklRcQm46V1uDpLodyJO6DiOLm3o5Se6Ano8uFuHOYmsy5CzsTzpuL74amCrIpLTc
R5cc7O2M3vpbvSQ54CZOn7mhpO8oAYWHkFtyi56CaTDXWm/+uYmxh3OU+PQhjJ98mxYbYLZIlioW
cfPW/Zr0H80GHSWNRP5QW6Qqt5Wv9jXbZxY3/carGpQOTpmKU287+Atnn6gAFosH5M1QVsWOOSgL
OvnG0232TNPSop8D9geqsQvXMUTpaaCi23H7qX2ZSJZVTulzIwkTxq+d81/XNp8u6U6MwOQMk2R2
9/HLkbI7/tr+98Wx31DAb4x+cC3LhFvD3/jxvDZfsQJHH8ZvwnrRPttWfFhJe21brcEkoxy5FQwG
+PFxzhPCTx7707jERE3xDO6SO+uCUCzkFAGhS9gBtgn5AATm2GMeqfPWiNwcbU67fCeDNUwLXtcX
PitKI+QkRSuBdhjza83K+uJl3Oax9v5CDEq7Tnqgda0KE4bqTE2HzusGQen02gcbikl6myK6+Yt4
qg9ap66q7oeXNWmzvlyriMRPW1jhlBDBs7+c8WXmaoEwp3/Q2/KOY1/iSWJ9me+98Xg8acVrowpl
yzak3DFmWl6pL1AOnUuyBwK9pcXv/Nd6YvZ5nvCHAML9b6lRL89CrQsJcPuyq+FARpFmNdK+rG8U
xSDsiNVMn/GU/p2fbsAliRSZvs6N4V/Rx2ou2NNH0dGxgyjjOiFxA07uzdlO6oTBRa3OwTbowIvu
1echlPdC81gpj1Y4qk3GF23GRNmg+szUHtgN3ZY6nkQyPi2jlzUnujxI18QjyrtljpkExv5npV6/
SYssfRGmk7+HJjx/Mut8mlg9ctOu06iMXN/FkxyQ6EA7LF/vqQfnoK6oZE9W4A+2n0G3C1uw+77V
bnfVTbZpjQ2QB//lTefrAo4ofuXOpnflZyLh9uw3/mOYAgrZdzNyQaSuSIyWZXiUK25I+fJ0KB4M
iPp3lTFB7T5QN+dj0sOsCV8h5Ddb1bGz3i3oXtWQA4BP0xBYU8I+A7XUnVT7lYUrcyqv/IZopU7K
RqUtg/qAnyvngyyAanWnSQ6FsozCWrTp9mUXsFRwVk5sRIQBplyXzCxN5Ard6mWp5l29zHz3xOkZ
YFoXavKtVC6IKVTwfHAznTTPh00rVBLizrERZxBCixRI6uKBZjRg75bpN9ZQdNntJLIu9oBpWEVh
mz9nDf9YsNAyWhTdis65M24WkS1TD16XNlia/VTa8x0KZSDhJQlO+DOdLf8lYDUzIQQWSqrObEjZ
ZUx7OG8hv0rmxPVST1PzyUeCAQpc9Gjx/uFJtuie3Hl0dYZcUOwRG0gx6WWKigR4Tghy8nkX2Vyn
YNod2CfiOahX8QkYUlmDOSBkZsX1T92ZV+62a344uUdP344ZRFfJBmUU/CZqhrdpwErn+0El47hW
uzYgW43iwBesIBEPXnBi
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity DVI_TX_Top is
port(
  I_rst_n :  in std_logic;
  I_serial_clk :  in std_logic;
  I_rgb_clk :  in std_logic;
  I_rgb_vs :  in std_logic;
  I_rgb_hs :  in std_logic;
  I_rgb_de :  in std_logic;
  I_rgb_r :  in std_logic_vector(7 downto 0);
  I_rgb_g :  in std_logic_vector(7 downto 0);
  I_rgb_b :  in std_logic_vector(7 downto 0);
  O_tmds_clk_p :  out std_logic;
  O_tmds_clk_n :  out std_logic;
  O_tmds_data_p :  out std_logic_vector(2 downto 0);
  O_tmds_data_n :  out std_logic_vector(2 downto 0));
end DVI_TX_Top;
architecture beh of DVI_TX_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~rgb2dvi.DVI_TX_Top\
port(
  I_rgb_clk: in std_logic;
  I_serial_clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  I_rst_n: in std_logic;
  I_rgb_de: in std_logic;
  I_rgb_vs: in std_logic;
  I_rgb_hs: in std_logic;
  I_rgb_r : in std_logic_vector(7 downto 0);
  I_rgb_g : in std_logic_vector(7 downto 0);
  I_rgb_b : in std_logic_vector(7 downto 0);
  O_tmds_clk_p: out std_logic;
  O_tmds_clk_n: out std_logic;
  O_tmds_data_p : out std_logic_vector(2 downto 0);
  O_tmds_data_n : out std_logic_vector(2 downto 0));
end component;
begin
GND_s3: GND
port map (
  G => GND_0);
VCC_s3: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
rgb2dvi_inst: \~rgb2dvi.DVI_TX_Top\
port map(
  I_rgb_clk => I_rgb_clk,
  I_serial_clk => I_serial_clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  I_rst_n => I_rst_n,
  I_rgb_de => I_rgb_de,
  I_rgb_vs => I_rgb_vs,
  I_rgb_hs => I_rgb_hs,
  I_rgb_r(7 downto 0) => I_rgb_r(7 downto 0),
  I_rgb_g(7 downto 0) => I_rgb_g(7 downto 0),
  I_rgb_b(7 downto 0) => I_rgb_b(7 downto 0),
  O_tmds_clk_p => O_tmds_clk_p,
  O_tmds_clk_n => O_tmds_clk_n,
  O_tmds_data_p(2 downto 0) => O_tmds_data_p(2 downto 0),
  O_tmds_data_n(2 downto 0) => O_tmds_data_n(2 downto 0));
end beh;
