library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- This contains 2.C of the AtoMMC2 firmware (10K x 16)

-- For f_log2 definition
use WORK.SynthCtrlPack.all;

entity XPM is
    generic (
        WIDTH : integer;
        SIZE  : integer
    );
    port(
        cp2     : in  std_logic;
        ce      : in  std_logic;
        address : in  std_logic_vector(f_log2(SIZE) - 1 downto 0);
        din     : in  std_logic_vector(WIDTH - 1 downto 0);
        dout    : out std_logic_vector(WIDTH - 1 downto 0);
        we      : in  std_logic
    );
end;

architecture RTL of XPM is
    
    type ram_type is array (0 to SIZE - 1) of std_logic_vector (WIDTH - 1 downto 0);

    signal RAM : ram_type := (
        x"940C",
        x"003D",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"0078",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"4F42",
        x"544F",
        x"5244",
        x"2E56",
        x"4643",
        x"0047",
        x"4F42",
        x"544F",
        x"5244",
        x"2E56",
        x"4643",
        x"0047",
        x"002A",
        x"2411",
        x"BE1F",
        x"EFCF",
        x"E0DF",
        x"BFDE",
        x"BFCD",
        x"E010",
        x"E6A0",
        x"E0B0",
        x"EBEE",
        x"E4F6",
        x"EF0F",
        x"9503",
        x"BF0B",
        x"C004",
        x"95D8",
        x"920D",
        x"9631",
        x"F3C8",
        x"39AE",
        x"07B1",
        x"F7C9",
        x"E01D",
        x"E9AE",
        x"E0B0",
        x"C001",
        x"921D",
        x"33A6",
        x"07B1",
        x"F7E1",
        x"940E",
        x"2211",
        x"940C",
        x"235D",
        x"940C",
        x"0000",
        x"9508",
        x"9508",
        x"CFFF",
        x"BA1A",
        x"B78A",
        x"7F8C",
        x"BF8A",
        x"B78A",
        x"6082",
        x"BF8A",
        x"B789",
        x"7F8C",
        x"BF89",
        x"98BC",
        x"9AC4",
        x"9AB8",
        x"9AC0",
        x"9AB9",
        x"9AC1",
        x"9ABB",
        x"98C3",
        x"988B",
        x"9508",
        x"921F",
        x"920F",
        x"B60F",
        x"920F",
        x"2411",
        x"900F",
        x"BE0F",
        x"900F",
        x"901F",
        x"9518",
        x"9A8B",
        x"9893",
        x"E98F",
        x"E09F",
        x"9701",
        x"F7F1",
        x"C000",
        x"0000",
        x"988B",
        x"9893",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"0F4E",
        x"1F5F",
        x"17E4",
        x"07F5",
        x"F039",
        x"9121",
        x"2FA8",
        x"2FB9",
        x"932D",
        x"2F8A",
        x"2F9B",
        x"CFF6",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F26",
        x"2F37",
        x"2FE6",
        x"2FF7",
        x"9639",
        x"2FA8",
        x"2FB9",
        x"961E",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9751",
        x"2B45",
        x"2B46",
        x"2B47",
        x"F409",
        x"C064",
        x"9652",
        x"91CD",
        x"91DC",
        x"9753",
        x"2F4C",
        x"2F5D",
        x"2F0E",
        x"2F1F",
        x"E080",
        x"E090",
        x"2FE0",
        x"2FF1",
        x"2FA4",
        x"2FB5",
        x"916D",
        x"2F4A",
        x"2F5B",
        x"3260",
        x"F081",
        x"3065",
        x"F409",
        x"EE65",
        x"2FE0",
        x"2FF1",
        x"9631",
        x"2FA0",
        x"2FB1",
        x"936C",
        x"9601",
        x"3088",
        x"0591",
        x"F019",
        x"2F0E",
        x"2F1F",
        x"CFE7",
        x"8588",
        x"3280",
        x"F119",
        x"E28E",
        x"2FAE",
        x"2FBF",
        x"938D",
        x"2EEA",
        x"2EFB",
        x"2F6C",
        x"2F7D",
        x"5F68",
        x"4F7F",
        x"2F8E",
        x"2F9F",
        x"9604",
        x"2DEE",
        x"2DFF",
        x"2FA6",
        x"2FB7",
        x"911D",
        x"2F6A",
        x"2F7B",
        x"3210",
        x"F069",
        x"2D4E",
        x"2D5F",
        x"5F4F",
        x"4F5F",
        x"8310",
        x"1748",
        x"0759",
        x"F019",
        x"2EE4",
        x"2EF5",
        x"CFEC",
        x"2FE8",
        x"2FF9",
        x"858B",
        x"2FA2",
        x"2FB3",
        x"9618",
        x"938C",
        x"9718",
        x"8D4C",
        x"8D5D",
        x"8D6E",
        x"8D7F",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9713",
        x"8D88",
        x"8D99",
        x"9615",
        x"939C",
        x"938E",
        x"9714",
        x"898E",
        x"899F",
        x"9617",
        x"939C",
        x"938E",
        x"9716",
        x"8210",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"22B6",
        x"E0A0",
        x"E0B0",
        x"E3E0",
        x"E0F1",
        x"940C",
        x"2294",
        x"2FC8",
        x"2FD9",
        x"2E84",
        x"2E95",
        x"2EA6",
        x"2EB7",
        x"A4CE",
        x"A4DF",
        x"A8E8",
        x"A8F9",
        x"16C4",
        x"06D5",
        x"06E6",
        x"06F7",
        x"F409",
        x"C052",
        x"818C",
        x"2388",
        x"F439",
        x"1481",
        x"0491",
        x"04A1",
        x"04B1",
        x"F409",
        x"C049",
        x"C038",
        x"A96A",
        x"A97B",
        x"E001",
        x"2D5F",
        x"2D4E",
        x"2D3D",
        x"2D2C",
        x"8189",
        x"940E",
        x"1809",
        x"2B89",
        x"F019",
        x"E081",
        x"E090",
        x"C03B",
        x"821C",
        x"8D8A",
        x"8D9B",
        x"8DAC",
        x"8DBD",
        x"A14A",
        x"A15B",
        x"A16C",
        x"A17D",
        x"0F84",
        x"1F95",
        x"1FA6",
        x"1FB7",
        x"16C8",
        x"06D9",
        x"06EA",
        x"06FB",
        x"F6C0",
        x"811B",
        x"3012",
        x"F2A8",
        x"8D8A",
        x"8D9B",
        x"8DAC",
        x"8DBD",
        x"0EC8",
        x"1ED9",
        x"1EEA",
        x"1EFB",
        x"A96A",
        x"A97B",
        x"E001",
        x"2D5F",
        x"2D4E",
        x"2D3D",
        x"2D2C",
        x"8189",
        x"940E",
        x"1809",
        x"5011",
        x"CFEA",
        x"A96A",
        x"A97B",
        x"E001",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"8189",
        x"940E",
        x"17FF",
        x"2B89",
        x"F641",
        x"A68E",
        x"A69F",
        x"AAA8",
        x"AAB9",
        x"E080",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"22B0",
        x"930F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"A98A",
        x"A99B",
        x"E001",
        x"2F24",
        x"2F35",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"8189",
        x"940E",
        x"17FF",
        x"2B89",
        x"F539",
        x"A9EA",
        x"A9FB",
        x"2FAE",
        x"2FBF",
        x"50A2",
        x"4FBE",
        x"918D",
        x"919C",
        x"3585",
        x"4A9A",
        x"F4C1",
        x"A986",
        x"A997",
        x"ADA0",
        x"ADB1",
        x"27BB",
        x"3486",
        x"4491",
        x"45A4",
        x"05B1",
        x"F081",
        x"5AEE",
        x"4FFF",
        x"8140",
        x"8151",
        x"8162",
        x"8173",
        x"2777",
        x"E081",
        x"3446",
        x"4451",
        x"4564",
        x"0571",
        x"F431",
        x"C002",
        x"E082",
        x"C003",
        x"E080",
        x"C001",
        x"E083",
        x"91DF",
        x"91CF",
        x"910F",
        x"9508",
        x"2FE8",
        x"2FF9",
        x"9700",
        x"F099",
        x"8180",
        x"2388",
        x"F081",
        x"8186",
        x"8197",
        x"1786",
        x"0797",
        x"F459",
        x"8181",
        x"940E",
        x"17FC",
        x"FF80",
        x"C003",
        x"E083",
        x"E090",
        x"9508",
        x"E080",
        x"E090",
        x"9508",
        x"E089",
        x"E090",
        x"9508",
        x"930F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"940E",
        x"012A",
        x"9700",
        x"F009",
        x"C06B",
        x"8188",
        x"3083",
        x"F009",
        x"C05A",
        x"818D",
        x"2388",
        x"F409",
        x"C056",
        x"A61E",
        x"A61F",
        x"AA18",
        x"AA19",
        x"A9EA",
        x"A9FB",
        x"2F8E",
        x"2F9F",
        x"5F9E",
        x"17E8",
        x"07F9",
        x"F011",
        x"9211",
        x"CFFB",
        x"A9EA",
        x"A9FB",
        x"2FAE",
        x"2FBF",
        x"50A2",
        x"4FBE",
        x"E585",
        x"EA9A",
        x"938D",
        x"939C",
        x"E582",
        x"E592",
        x"E6A1",
        x"E4B1",
        x"8380",
        x"8391",
        x"83A2",
        x"83B3",
        x"2F2E",
        x"2F3F",
        x"512C",
        x"4F3E",
        x"E742",
        x"E752",
        x"E461",
        x"E671",
        x"2FA2",
        x"2FB3",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9713",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"2F2E",
        x"2F3F",
        x"5128",
        x"4F3E",
        x"2FA2",
        x"2FB3",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9713",
        x"854A",
        x"855B",
        x"856C",
        x"857D",
        x"2FAE",
        x"2FBF",
        x"51A4",
        x"4FBE",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9713",
        x"892A",
        x"893B",
        x"894C",
        x"895D",
        x"E001",
        x"2F6E",
        x"2F7F",
        x"8189",
        x"940E",
        x"1809",
        x"821D",
        x"E040",
        x"E050",
        x"E060",
        x"8189",
        x"940E",
        x"1813",
        x"E031",
        x"E020",
        x"2B89",
        x"F409",
        x"E030",
        x"2F83",
        x"2F92",
        x"91DF",
        x"91CF",
        x"910F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E7E5",
        x"E0F2",
        x"940C",
        x"2293",
        x"2FC8",
        x"2FD9",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"C0A8",
        x"8D8E",
        x"8D9F",
        x"A1A8",
        x"A1B9",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C09E",
        x"A08A",
        x"A09B",
        x"A0AC",
        x"A0BD",
        x"8188",
        x"3082",
        x"F409",
        x"C051",
        x"3083",
        x"F409",
        x"C06B",
        x"3081",
        x"F009",
        x"C08B",
        x"2F04",
        x"2F15",
        x"9516",
        x"9507",
        x"0D0C",
        x"1D1D",
        x"2F80",
        x"2F91",
        x"2F89",
        x"2799",
        x"9586",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"012A",
        x"2B89",
        x"F009",
        x"C071",
        x"2F80",
        x"2F91",
        x"7091",
        x"A9EA",
        x"A9FB",
        x"0FE8",
        x"1FF9",
        x"8070",
        x"5F0F",
        x"4F1F",
        x"2F80",
        x"2F91",
        x"2F89",
        x"2799",
        x"9586",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"012A",
        x"2B89",
        x"F009",
        x"C053",
        x"7011",
        x"A9EA",
        x"A9FB",
        x"0FE0",
        x"1FF1",
        x"8180",
        x"2D67",
        x"E070",
        x"2B78",
        x"FEC0",
        x"C006",
        x"E044",
        x"9576",
        x"9567",
        x"954A",
        x"F7E1",
        x"C01C",
        x"707F",
        x"C01A",
        x"2F45",
        x"2F56",
        x"2F67",
        x"2777",
        x"0D48",
        x"1D59",
        x"1D6A",
        x"1D7B",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"012A",
        x"2B89",
        x"F591",
        x"0CCC",
        x"1CDD",
        x"94E8",
        x"F8C0",
        x"E081",
        x"22D8",
        x"A9EA",
        x"A9FB",
        x"0DEC",
        x"1DFD",
        x"8160",
        x"8171",
        x"E080",
        x"E090",
        x"C02C",
        x"E097",
        x"9576",
        x"9567",
        x"9557",
        x"9547",
        x"959A",
        x"F7D1",
        x"0D48",
        x"1D59",
        x"1D6A",
        x"1D7B",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"012A",
        x"2B89",
        x"F491",
        x"0CCC",
        x"1CDD",
        x"0CCC",
        x"1CDD",
        x"EF8C",
        x"22C8",
        x"E081",
        x"22D8",
        x"A9EA",
        x"A9FB",
        x"0DEC",
        x"1DFD",
        x"8160",
        x"8171",
        x"8182",
        x"8193",
        x"709F",
        x"C009",
        x"EF6F",
        x"EF7F",
        x"EF8F",
        x"EF9F",
        x"C004",
        x"E061",
        x"E070",
        x"E080",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0ED",
        x"940C",
        x"22AF",
        x"E0A8",
        x"E0B0",
        x"E3E8",
        x"E0F3",
        x"940C",
        x"2290",
        x"2E88",
        x"2E99",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"8309",
        x"831A",
        x"832B",
        x"833C",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"C0F0",
        x"2FE8",
        x"2FF9",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C0E4",
        x"A042",
        x"A053",
        x"A064",
        x"A075",
        x"8180",
        x"3082",
        x"F409",
        x"C088",
        x"3083",
        x"F409",
        x"C0A7",
        x"3081",
        x"F009",
        x"C0CE",
        x"2EA4",
        x"2EB5",
        x"94B6",
        x"94A7",
        x"0CAC",
        x"1CBD",
        x"2D8A",
        x"2D9B",
        x"2F89",
        x"2799",
        x"9586",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2D88",
        x"2D99",
        x"940E",
        x"012A",
        x"9700",
        x"F009",
        x"C0B6",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"912D",
        x"913C",
        x"97D3",
        x"2D8A",
        x"2D9B",
        x"7091",
        x"0F28",
        x"1F39",
        x"2DBF",
        x"2DAE",
        x"2D9D",
        x"2D8C",
        x"7081",
        x"2799",
        x"27AA",
        x"27BB",
        x"838D",
        x"839E",
        x"83AF",
        x"87B8",
        x"FEC0",
        x"C009",
        x"2FA2",
        x"2FB3",
        x"919C",
        x"709F",
        x"8189",
        x"9582",
        x"7F80",
        x"2B89",
        x"C001",
        x"8189",
        x"2FE2",
        x"2FF3",
        x"8380",
        x"EFFF",
        x"1AAF",
        x"0ABF",
        x"E081",
        x"2DA8",
        x"2DB9",
        x"9614",
        x"938C",
        x"2D8A",
        x"2D9B",
        x"2F89",
        x"2799",
        x"9586",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2D88",
        x"2D99",
        x"940E",
        x"012A",
        x"9700",
        x"F009",
        x"C074",
        x"E0B1",
        x"22BB",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"0DEA",
        x"1DFB",
        x"812D",
        x"813E",
        x"814F",
        x"8558",
        x"2B23",
        x"2B24",
        x"2B25",
        x"F069",
        x"8049",
        x"805A",
        x"806B",
        x"807C",
        x"E024",
        x"9476",
        x"9467",
        x"9457",
        x"9447",
        x"952A",
        x"F7D1",
        x"2D24",
        x"C005",
        x"8120",
        x"7F20",
        x"813A",
        x"703F",
        x"2B23",
        x"8320",
        x"C04E",
        x"2F45",
        x"2F56",
        x"2F67",
        x"2777",
        x"0D44",
        x"1D55",
        x"1D66",
        x"1D77",
        x"2D88",
        x"2D99",
        x"940E",
        x"012A",
        x"9700",
        x"F009",
        x"C03F",
        x"0CCC",
        x"1CDD",
        x"94E8",
        x"F8C0",
        x"E031",
        x"22D3",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"0DEC",
        x"1DFD",
        x"8129",
        x"813A",
        x"8331",
        x"8320",
        x"C02C",
        x"E0F7",
        x"9576",
        x"9567",
        x"9557",
        x"9547",
        x"95FA",
        x"F7D1",
        x"0D44",
        x"1D55",
        x"1D66",
        x"1D77",
        x"2D88",
        x"2D99",
        x"940E",
        x"012A",
        x"9700",
        x"F4D9",
        x"0CCC",
        x"1CDD",
        x"0CCC",
        x"1CDD",
        x"EF3C",
        x"22C3",
        x"E031",
        x"22D3",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"0DEC",
        x"1DFD",
        x"8129",
        x"813A",
        x"814B",
        x"815C",
        x"8320",
        x"8331",
        x"8342",
        x"8353",
        x"C002",
        x"E082",
        x"E090",
        x"E021",
        x"2DA8",
        x"2DB9",
        x"9614",
        x"932C",
        x"C002",
        x"E082",
        x"E090",
        x"9628",
        x"E1E0",
        x"940C",
        x"22AC",
        x"E0A4",
        x"E0B0",
        x"E4E4",
        x"E0F4",
        x"940C",
        x"228E",
        x"2E28",
        x"2E39",
        x"2E44",
        x"2E55",
        x"2E66",
        x"2E77",
        x"2FA8",
        x"2FB9",
        x"965E",
        x"912D",
        x"913D",
        x"914D",
        x"915C",
        x"9791",
        x"8329",
        x"833A",
        x"834B",
        x"835C",
        x"1441",
        x"0451",
        x"0461",
        x"0471",
        x"F489",
        x"961A",
        x"908D",
        x"909D",
        x"90AD",
        x"90BC",
        x"971D",
        x"1481",
        x"0491",
        x"04A1",
        x"04B1",
        x"F111",
        x"1682",
        x"0693",
        x"06A4",
        x"06B5",
        x"F4E8",
        x"C021",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"940E",
        x"026F",
        x"3062",
        x"0571",
        x"0581",
        x"0591",
        x"F410",
        x"E041",
        x"C02D",
        x"8129",
        x"813A",
        x"814B",
        x"815C",
        x"1762",
        x"0773",
        x"0784",
        x"0795",
        x"F408",
        x"C09A",
        x"2CB7",
        x"2CA6",
        x"2C95",
        x"2C84",
        x"C005",
        x"2488",
        x"9483",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"2CFB",
        x"2CEA",
        x"2CD9",
        x"2CC8",
        x"EF3F",
        x"1AC3",
        x"0AD3",
        x"0AE3",
        x"0AF3",
        x"8129",
        x"813A",
        x"814B",
        x"815C",
        x"16C2",
        x"06D3",
        x"06E4",
        x"06F5",
        x"F080",
        x"E032",
        x"1683",
        x"0491",
        x"04A1",
        x"04B1",
        x"F428",
        x"E040",
        x"E030",
        x"E020",
        x"E090",
        x"C076",
        x"E062",
        x"2EC6",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2D82",
        x"2D93",
        x"940E",
        x"026F",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F0C1",
        x"3F6F",
        x"EF4F",
        x"0774",
        x"0784",
        x"0794",
        x"F429",
        x"EF4F",
        x"EF3F",
        x"EF2F",
        x"EF9F",
        x"C059",
        x"3061",
        x"0571",
        x"0581",
        x"0591",
        x"F409",
        x"CFAA",
        x"14C8",
        x"04D9",
        x"04EA",
        x"04FB",
        x"F009",
        x"CFBE",
        x"CFD1",
        x"EF0F",
        x"EF1F",
        x"EF2F",
        x"E03F",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2D82",
        x"2D93",
        x"940E",
        x"0332",
        x"2B89",
        x"F701",
        x"1441",
        x"0451",
        x"0461",
        x"0471",
        x"F509",
        x"2DA2",
        x"2DB3",
        x"961A",
        x"92CD",
        x"92DD",
        x"92ED",
        x"92FC",
        x"971D",
        x"961E",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9751",
        x"3F4F",
        x"EFBF",
        x"075B",
        x"076B",
        x"077B",
        x"F0E9",
        x"5041",
        x"0951",
        x"0961",
        x"0971",
        x"2DE2",
        x"2DF3",
        x"8746",
        x"8757",
        x"8B60",
        x"8B71",
        x"E081",
        x"8385",
        x"C010",
        x"2D3F",
        x"2D2E",
        x"2D1D",
        x"2D0C",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"2D82",
        x"2D93",
        x"940E",
        x"0332",
        x"2B89",
        x"F009",
        x"CFAB",
        x"CFCF",
        x"2D4C",
        x"2D3D",
        x"2D2E",
        x"2D9F",
        x"C003",
        x"2F46",
        x"2F37",
        x"2F28",
        x"2F64",
        x"2F73",
        x"2F82",
        x"9624",
        x"E1E2",
        x"940C",
        x"22AA",
        x"E0A0",
        x"E0B0",
        x"E2ED",
        x"E0F5",
        x"940C",
        x"2293",
        x"2FC8",
        x"2FD9",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"C05E",
        x"8D8E",
        x"8D9F",
        x"A1A8",
        x"A1B9",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C054",
        x"2477",
        x"9473",
        x"8D8E",
        x"8D9F",
        x"A1A8",
        x"A1B9",
        x"16C8",
        x"06D9",
        x"06EA",
        x"06FB",
        x"F488",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"026F",
        x"2E86",
        x"2E97",
        x"2EA8",
        x"2EB9",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F419",
        x"E080",
        x"E090",
        x"C037",
        x"E081",
        x"1688",
        x"0491",
        x"04A1",
        x"04B1",
        x"F179",
        x"EF8F",
        x"1688",
        x"0698",
        x"06A8",
        x"06B8",
        x"F131",
        x"E000",
        x"E010",
        x"E020",
        x"E030",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"0332",
        x"9700",
        x"F4E9",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"3F4F",
        x"EF8F",
        x"0758",
        x"0768",
        x"0778",
        x"F049",
        x"5F4F",
        x"4F5F",
        x"4F6F",
        x"4F7F",
        x"874E",
        x"875F",
        x"8B68",
        x"8B79",
        x"827D",
        x"2CFB",
        x"2CEA",
        x"2CD9",
        x"2CC8",
        x"CFB1",
        x"E081",
        x"E090",
        x"C002",
        x"E082",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0ED",
        x"940C",
        x"22AF",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"5042",
        x"0951",
        x"0961",
        x"0971",
        x"8D8E",
        x"8D9F",
        x"A1A8",
        x"A1B9",
        x"9702",
        x"09A1",
        x"09B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F4D8",
        x"80CA",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"2F97",
        x"2F86",
        x"2F75",
        x"2F64",
        x"2D5F",
        x"2D4E",
        x"2D3D",
        x"2D2C",
        x"940E",
        x"226A",
        x"2E82",
        x"2E93",
        x"2EA4",
        x"2EB5",
        x"A56A",
        x"A57B",
        x"A58C",
        x"A59D",
        x"0D68",
        x"1D79",
        x"1D8A",
        x"1D9B",
        x"C004",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F06",
        x"2F17",
        x"837D",
        x"836C",
        x"814E",
        x"815F",
        x"8568",
        x"8579",
        x"3041",
        x"0551",
        x"0561",
        x"0571",
        x"F419",
        x"E082",
        x"E090",
        x"C08F",
        x"81E8",
        x"81F9",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F790",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F549",
        x"8180",
        x"3083",
        x"F449",
        x"A146",
        x"A157",
        x"A560",
        x"A571",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F4E9",
        x"861A",
        x"861B",
        x"861C",
        x"861D",
        x"8580",
        x"8591",
        x"1708",
        x"0719",
        x"F6C0",
        x"A186",
        x"A197",
        x"A5A0",
        x"A5B1",
        x"2F20",
        x"2F31",
        x"E044",
        x"9536",
        x"9527",
        x"954A",
        x"F7E1",
        x"0F82",
        x"1F93",
        x"1DA1",
        x"1DB1",
        x"878E",
        x"879F",
        x"8BA8",
        x"8BB9",
        x"C042",
        x"80E2",
        x"2CF1",
        x"E084",
        x"0CEE",
        x"1CFF",
        x"958A",
        x"F7E1",
        x"8188",
        x"8199",
        x"150E",
        x"051F",
        x"F108",
        x"940E",
        x"026F",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"3F4F",
        x"EF8F",
        x"0758",
        x"0768",
        x"0778",
        x"F1E1",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"CFA6",
        x"81E8",
        x"81F9",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"CF9A",
        x"190E",
        x"091F",
        x"CFDA",
        x"874A",
        x"875B",
        x"876C",
        x"877D",
        x"940E",
        x"059E",
        x"2F20",
        x"2F31",
        x"E0B4",
        x"9536",
        x"9527",
        x"95BA",
        x"F7E1",
        x"0F62",
        x"1F73",
        x"1D81",
        x"1D91",
        x"876E",
        x"877F",
        x"8B88",
        x"8B99",
        x"81E8",
        x"81F9",
        x"700F",
        x"2711",
        x"E0A5",
        x"0F00",
        x"1F11",
        x"95AA",
        x"F7E1",
        x"A982",
        x"A993",
        x"0F80",
        x"1F91",
        x"8B9B",
        x"8B8A",
        x"E080",
        x"E090",
        x"C002",
        x"E081",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"22B6",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"816C",
        x"817D",
        x"940E",
        x"05E4",
        x"9700",
        x"F491",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"9700",
        x"F441",
        x"89EA",
        x"89FB",
        x"EE25",
        x"8320",
        x"81E8",
        x"81F9",
        x"E021",
        x"8324",
        x"91DF",
        x"91CF",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"EBE5",
        x"E0F6",
        x"940C",
        x"2294",
        x"2FC8",
        x"2FD9",
        x"2EC6",
        x"2ED7",
        x"810C",
        x"811D",
        x"5F0F",
        x"4F1F",
        x"1501",
        x"0511",
        x"F419",
        x"E084",
        x"E090",
        x"C0F9",
        x"858E",
        x"859F",
        x"89A8",
        x"89B9",
        x"9700",
        x"05A1",
        x"05B1",
        x"F3A9",
        x"2EE0",
        x"2EF1",
        x"E02F",
        x"22E2",
        x"24FF",
        x"14E1",
        x"04F1",
        x"F009",
        x"C0D4",
        x"9601",
        x"1DA1",
        x"1DB1",
        x"878E",
        x"879F",
        x"8BA8",
        x"8BB9",
        x"854A",
        x"855B",
        x"856C",
        x"857D",
        x"8188",
        x"8199",
        x"2FE8",
        x"2FF9",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F431",
        x"8580",
        x"8591",
        x"1708",
        x"0719",
        x"F698",
        x"C0BA",
        x"8122",
        x"E030",
        x"5021",
        x"0931",
        x"2FE0",
        x"2FF1",
        x"E0A4",
        x"95F6",
        x"95E7",
        x"95AA",
        x"F7E1",
        x"232E",
        x"233F",
        x"2B23",
        x"F009",
        x"C0AA",
        x"940E",
        x"026F",
        x"2E86",
        x"2E97",
        x"2EA8",
        x"2EB9",
        x"3062",
        x"0571",
        x"0581",
        x"0591",
        x"F418",
        x"E082",
        x"E090",
        x"C0B0",
        x"3F6F",
        x"EF2F",
        x"0772",
        x"0782",
        x"0792",
        x"F419",
        x"E081",
        x"E090",
        x"C0A7",
        x"8188",
        x"8199",
        x"2FE8",
        x"2FF9",
        x"8D46",
        x"8D57",
        x"A160",
        x"A171",
        x"1684",
        x"0695",
        x"06A6",
        x"06B7",
        x"F408",
        x"C075",
        x"14C1",
        x"04D1",
        x"F409",
        x"CF99",
        x"854A",
        x"855B",
        x"856C",
        x"857D",
        x"940E",
        x"043E",
        x"2E86",
        x"2E97",
        x"2EA8",
        x"2EB9",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F409",
        x"C083",
        x"3061",
        x"0571",
        x"0581",
        x"0591",
        x"F269",
        x"3F6F",
        x"EF2F",
        x"0772",
        x"0782",
        x"0792",
        x"F281",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"2B89",
        x"F631",
        x"81E8",
        x"81F9",
        x"A802",
        x"A9F3",
        x"2DE0",
        x"2F8E",
        x"2F9F",
        x"5F9E",
        x"17E8",
        x"07F9",
        x"F011",
        x"9211",
        x"CFFB",
        x"80C8",
        x"80D9",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"059E",
        x"2DEC",
        x"2DFD",
        x"A766",
        x"A777",
        x"AB80",
        x"AB91",
        x"2CD1",
        x"24CC",
        x"94C3",
        x"81E8",
        x"81F9",
        x"8182",
        x"16D8",
        x"F4D8",
        x"82C4",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"2B89",
        x"F009",
        x"CF95",
        x"81E8",
        x"81F9",
        x"A586",
        x"A597",
        x"A9A0",
        x"A9B1",
        x"9601",
        x"1DA1",
        x"1DB1",
        x"A786",
        x"A797",
        x"ABA0",
        x"ABB1",
        x"94D3",
        x"CFE0",
        x"A586",
        x"A597",
        x"A9A0",
        x"A9B1",
        x"198D",
        x"0991",
        x"09A1",
        x"09B1",
        x"A786",
        x"A797",
        x"ABA0",
        x"ABB1",
        x"868A",
        x"869B",
        x"86AC",
        x"86BD",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"8188",
        x"8199",
        x"940E",
        x"059E",
        x"876E",
        x"877F",
        x"8B88",
        x"8B99",
        x"831D",
        x"830C",
        x"81E8",
        x"81F9",
        x"E055",
        x"0CEE",
        x"1CFF",
        x"955A",
        x"F7E1",
        x"A982",
        x"A993",
        x"0D8E",
        x"1D9F",
        x"8B9B",
        x"8B8A",
        x"E080",
        x"E090",
        x"C002",
        x"E087",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"22B0",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"927F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F06",
        x"2F17",
        x"2FA6",
        x"2FB7",
        x"918C",
        x"5F6F",
        x"4F7F",
        x"3280",
        x"F3B9",
        x"328F",
        x"F011",
        x"358C",
        x"F439",
        x"5F0F",
        x"4F1F",
        x"821E",
        x"821F",
        x"8618",
        x"8619",
        x"C00A",
        x"81E8",
        x"81F9",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"838E",
        x"839F",
        x"87A8",
        x"87B9",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"3280",
        x"F448",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"05E4",
        x"8A1B",
        x"8A1A",
        x"C113",
        x"E2B0",
        x"2EAB",
        x"E085",
        x"2EB8",
        x"89EC",
        x"89FD",
        x"2F8E",
        x"2F9F",
        x"960B",
        x"2FAE",
        x"2FBF",
        x"17A8",
        x"07B9",
        x"F011",
        x"92AD",
        x"CFFB",
        x"2FA0",
        x"2FB1",
        x"918C",
        x"328E",
        x"F051",
        x"2E20",
        x"2E31",
        x"E080",
        x"E090",
        x"E040",
        x"E050",
        x"E028",
        x"E030",
        x"2C91",
        x"C038",
        x"2F20",
        x"2F31",
        x"2F6E",
        x"2F7F",
        x"E080",
        x"E090",
        x"9601",
        x"2FA2",
        x"2FB3",
        x"914D",
        x"2F2A",
        x"2F3B",
        x"324E",
        x"F451",
        x"3083",
        x"0591",
        x"F409",
        x"C0E0",
        x"2FA6",
        x"2FB7",
        x"934D",
        x"2F6A",
        x"2F7B",
        x"CFEE",
        x"324F",
        x"F029",
        x"354C",
        x"F019",
        x"3241",
        x"F008",
        x"C0D3",
        x"0F08",
        x"1F19",
        x"3241",
        x"F410",
        x"E284",
        x"C001",
        x"E280",
        x"8783",
        x"C06D",
        x"327F",
        x"F1A9",
        x"357C",
        x"F199",
        x"327E",
        x"F4A9",
        x"3028",
        x"0531",
        x"F009",
        x"C0C0",
        x"0C99",
        x"0C99",
        x"E088",
        x"E090",
        x"E02B",
        x"E030",
        x"5F4F",
        x"4F5F",
        x"2DA2",
        x"2DB3",
        x"917D",
        x"2E2A",
        x"2E3B",
        x"2E77",
        x"3271",
        x"F730",
        x"C01A",
        x"1782",
        x"0793",
        x"F00C",
        x"C0AB",
        x"FD77",
        x"C0A9",
        x"2EE7",
        x"2CF1",
        x"E9A3",
        x"2E4A",
        x"E0A0",
        x"2E5A",
        x"2DA4",
        x"2DB5",
        x"90CD",
        x"2E4A",
        x"2E5B",
        x"20CC",
        x"F121",
        x"24DD",
        x"FCC7",
        x"94D0",
        x"14CE",
        x"04DF",
        x"F799",
        x"C095",
        x"E064",
        x"C001",
        x"E060",
        x"2B89",
        x"F409",
        x"C08F",
        x"8180",
        x"3E85",
        x"F409",
        x"82B0",
        x"3028",
        x"0531",
        x"F411",
        x"0C99",
        x"0C99",
        x"2D89",
        x"7083",
        x"3081",
        x"F409",
        x"6160",
        x"2D89",
        x"708C",
        x"3084",
        x"F409",
        x"6068",
        x"0F04",
        x"1F15",
        x"8763",
        x"C01B",
        x"EB6F",
        x"0F67",
        x"316A",
        x"F420",
        x"2DB9",
        x"60B2",
        x"2E9B",
        x"C00A",
        x"E96F",
        x"0F67",
        x"316A",
        x"F430",
        x"2D69",
        x"6061",
        x"2E96",
        x"EE60",
        x"2E76",
        x"0E77",
        x"2F6E",
        x"2F7F",
        x"0F68",
        x"1F79",
        x"2FA6",
        x"2FB7",
        x"927C",
        x"9601",
        x"CFA3",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"05E4",
        x"9700",
        x"F551",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"9700",
        x"F501",
        x"89EA",
        x"89FB",
        x"8180",
        x"2388",
        x"F0B1",
        x"8583",
        x"FD83",
        x"C00C",
        x"89AC",
        x"89BD",
        x"2F8E",
        x"2F9F",
        x"960B",
        x"17E8",
        x"07F9",
        x"F071",
        x"9131",
        x"912D",
        x"1732",
        x"F3C9",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"06AF",
        x"CFD9",
        x"E084",
        x"E090",
        x"C002",
        x"E080",
        x"E090",
        x"89EC",
        x"89FD",
        x"8523",
        x"7024",
        x"9700",
        x"F031",
        x"3084",
        x"0591",
        x"F521",
        x"2322",
        x"F0E9",
        x"C021",
        x"2322",
        x"F4F9",
        x"89EA",
        x"89FB",
        x"8583",
        x"FF84",
        x"C015",
        x"8984",
        x"8995",
        x"E0A0",
        x"E0B0",
        x"2FA8",
        x"2FB9",
        x"2799",
        x"2788",
        x"8D42",
        x"8D53",
        x"E060",
        x"E070",
        x"2B84",
        x"2B95",
        x"2BA6",
        x"2BB7",
        x"838E",
        x"839F",
        x"87A8",
        x"87B9",
        x"CEF6",
        x"E085",
        x"E090",
        x"C002",
        x"E086",
        x"E090",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"907F",
        x"905F",
        x"904F",
        x"903F",
        x"902F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"E060",
        x"E070",
        x"940E",
        x"05E4",
        x"2F08",
        x"2F19",
        x"9700",
        x"F009",
        x"C045",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"2F08",
        x"2F19",
        x"9700",
        x"F5C9",
        x"89EA",
        x"89FB",
        x"8180",
        x"3E85",
        x"F049",
        x"2388",
        x"F039",
        x"E061",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"06AF",
        x"CFE1",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"2F08",
        x"2F19",
        x"9700",
        x"F4F9",
        x"88EA",
        x"88FB",
        x"2DEE",
        x"2DFF",
        x"2D8E",
        x"2D9F",
        x"9680",
        x"17E8",
        x"07F9",
        x"F011",
        x"9211",
        x"CFFB",
        x"896C",
        x"897D",
        x"E04B",
        x"E050",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"0099",
        x"89EC",
        x"89FD",
        x"8583",
        x"7188",
        x"2DEE",
        x"2DFF",
        x"8784",
        x"81E8",
        x"81F9",
        x"E081",
        x"8384",
        x"2F80",
        x"2F91",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"22B6",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"E024",
        x"E030",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F0D9",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"9700",
        x"F519",
        x"89EA",
        x"89FB",
        x"8120",
        x"2322",
        x"F0E1",
        x"3E25",
        x"F019",
        x"8523",
        x"FF23",
        x"C01C",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"06AF",
        x"9700",
        x"F489",
        x"E020",
        x"E030",
        x"CFDC",
        x"2F82",
        x"2F93",
        x"1521",
        x"0531",
        x"F061",
        x"861E",
        x"861F",
        x"8A18",
        x"8A19",
        x"2F82",
        x"2F93",
        x"C005",
        x"E084",
        x"E090",
        x"2F28",
        x"2F39",
        x"CFF4",
        x"91DF",
        x"91CF",
        x"9508",
        x"2F68",
        x"2F79",
        x"EA88",
        x"E093",
        x"940E",
        x"00A8",
        x"9508",
        x"E0A8",
        x"E0B0",
        x"ECEB",
        x"E0F9",
        x"940C",
        x"2290",
        x"2F14",
        x"2FA8",
        x"2FB9",
        x"91ED",
        x"91FC",
        x"9711",
        x"8120",
        x"2733",
        x"FD27",
        x"9530",
        x"5320",
        x"0931",
        x"302A",
        x"0531",
        x"F438",
        x"8141",
        x"334A",
        x"F421",
        x"9632",
        x"93ED",
        x"93FC",
        x"C003",
        x"9120",
        x"009E",
        x"E030",
        x"2B23",
        x"F009",
        x"C107",
        x"9080",
        x"00A1",
        x"9090",
        x"00A2",
        x"2FE6",
        x"2FF7",
        x"8291",
        x"8280",
        x"1481",
        x"0491",
        x"F409",
        x"C0FE",
        x"2DA8",
        x"2DB9",
        x"918C",
        x"2388",
        x"F061",
        x"9611",
        x"918C",
        x"940E",
        x"17FC",
        x"FD80",
        x"C006",
        x"2311",
        x"F409",
        x"C13D",
        x"FD82",
        x"C141",
        x"C13A",
        x"2DE8",
        x"2DF9",
        x"8210",
        x"8211",
        x"E080",
        x"940E",
        x"17F9",
        x"FD80",
        x"C134",
        x"2311",
        x"F011",
        x"FD82",
        x"C133",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2D88",
        x"2D99",
        x"940E",
        x"0199",
        x"3081",
        x"F509",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"918D",
        x"919C",
        x"97D3",
        x"2FE8",
        x"2FF9",
        x"53EE",
        x"4FFE",
        x"8120",
        x"2322",
        x"F419",
        x"E08D",
        x"E090",
        x"C191",
        x"2FE8",
        x"2FF9",
        x"53EA",
        x"4FFE",
        x"8040",
        x"8051",
        x"8062",
        x"8073",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"2D88",
        x"2D99",
        x"940E",
        x"0199",
        x"C004",
        x"2C41",
        x"2C51",
        x"2C61",
        x"2C71",
        x"3083",
        x"F409",
        x"C104",
        x"2388",
        x"F719",
        x"2DE8",
        x"2DF9",
        x"A8A2",
        x"A8B3",
        x"2DAA",
        x"2DBB",
        x"961B",
        x"918D",
        x"919C",
        x"971C",
        x"1581",
        x"4092",
        x"F6B1",
        x"2DEA",
        x"2DFB",
        x"8966",
        x"8977",
        x"E080",
        x"E090",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F421",
        x"A164",
        x"A175",
        x"A186",
        x"A197",
        x"2DA8",
        x"2DB9",
        x"965A",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"975D",
        x"2DEA",
        x"2DFB",
        x"8920",
        x"9613",
        x"932C",
        x"E030",
        x"E040",
        x"E050",
        x"940E",
        x"226A",
        x"2EC2",
        x"2ED3",
        x"2EE4",
        x"2EF5",
        x"2DAA",
        x"2DBB",
        x"961E",
        x"918D",
        x"919C",
        x"971F",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"0F28",
        x"1F39",
        x"1D41",
        x"1D51",
        x"8329",
        x"833A",
        x"834B",
        x"835C",
        x"2DA8",
        x"2DB9",
        x"9692",
        x"932D",
        x"933D",
        x"934D",
        x"935C",
        x"9795",
        x"2DEA",
        x"2DFB",
        x"8515",
        x"9612",
        x"931C",
        x"9712",
        x"8921",
        x"8932",
        x"9619",
        x"933C",
        x"932E",
        x"9718",
        x"8983",
        x"8994",
        x"E0A0",
        x"E0B0",
        x"9700",
        x"05A1",
        x"05B1",
        x"F421",
        x"A180",
        x"A191",
        x"A1A2",
        x"A1B3",
        x"E044",
        x"9536",
        x"9527",
        x"954A",
        x"F7E1",
        x"2F42",
        x"2F53",
        x"E060",
        x"E070",
        x"834D",
        x"835E",
        x"836F",
        x"8778",
        x"2DEA",
        x"2DFB",
        x"8526",
        x"8537",
        x"2F68",
        x"2F79",
        x"2F8A",
        x"2F9B",
        x"1B62",
        x"0B73",
        x"0981",
        x"0991",
        x"196C",
        x"097D",
        x"098E",
        x"099F",
        x"812D",
        x"813E",
        x"814F",
        x"8558",
        x"1B62",
        x"0B73",
        x"0B84",
        x"0B95",
        x"2F21",
        x"E030",
        x"E040",
        x"E050",
        x"940E",
        x"2241",
        x"5F2E",
        x"4F3F",
        x"4F4F",
        x"4F5F",
        x"2DA8",
        x"2DB9",
        x"965E",
        x"932D",
        x"933D",
        x"934D",
        x"935C",
        x"9791",
        x"3F27",
        x"E0BF",
        x"073B",
        x"0541",
        x"0551",
        x"F408",
        x"C0C5",
        x"3F27",
        x"4F3F",
        x"0541",
        x"0551",
        x"F440",
        x"E012",
        x"C0BF",
        x"E08B",
        x"E090",
        x"C0CB",
        x"E08C",
        x"E090",
        x"C0C8",
        x"2DEA",
        x"2DFB",
        x"A584",
        x"A595",
        x"A5A6",
        x"A5B7",
        x"2DE8",
        x"2DF9",
        x"A386",
        x"A397",
        x"A7A0",
        x"A7B1",
        x"E013",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"812D",
        x"813E",
        x"814F",
        x"8558",
        x"0F82",
        x"1F93",
        x"1FA4",
        x"1FB5",
        x"0D8C",
        x"1D9D",
        x"1DAE",
        x"1DBF",
        x"2DE8",
        x"2DF9",
        x"A782",
        x"A793",
        x"A7A4",
        x"A7B5",
        x"EF8F",
        x"EF9F",
        x"EFAF",
        x"EFBF",
        x"8786",
        x"8797",
        x"8BA0",
        x"8BB1",
        x"8214",
        x"3013",
        x"F141",
        x"2DA8",
        x"2DB9",
        x"931C",
        x"2DE8",
        x"2DF9",
        x"A616",
        x"A617",
        x"AA10",
        x"AA11",
        x"9656",
        x"921D",
        x"921D",
        x"921D",
        x"921C",
        x"9759",
        x"9180",
        x"009F",
        x"9190",
        x"00A0",
        x"9601",
        x"9390",
        x"00A0",
        x"9380",
        x"009F",
        x"9617",
        x"939C",
        x"938E",
        x"9716",
        x"E080",
        x"E090",
        x"C07B",
        x"E083",
        x"E090",
        x"C078",
        x"E08A",
        x"E090",
        x"C075",
        x"E081",
        x"E090",
        x"C072",
        x"8215",
        x"2DAA",
        x"2DBB",
        x"96D0",
        x"918D",
        x"919C",
        x"97D1",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"0F28",
        x"1F39",
        x"1D41",
        x"1D51",
        x"8B22",
        x"8B33",
        x"8B44",
        x"8B55",
        x"E001",
        x"2D6A",
        x"2D7B",
        x"8181",
        x"940E",
        x"17FF",
        x"2B89",
        x"F009",
        x"CFBC",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"2FAE",
        x"2FBF",
        x"50A2",
        x"4FBE",
        x"918D",
        x"919C",
        x"3585",
        x"4A9A",
        x"F009",
        x"CFAC",
        x"8180",
        x"8191",
        x"81A2",
        x"81B3",
        x"3582",
        x"4592",
        x"46A1",
        x"44B1",
        x"F009",
        x"CFA2",
        x"2FAE",
        x"2FBF",
        x"51AC",
        x"4FBE",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"3782",
        x"4792",
        x"44A1",
        x"46B1",
        x"F009",
        x"CF93",
        x"2FAE",
        x"2FBF",
        x"51A4",
        x"4FBE",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"2DA8",
        x"2DB9",
        x"961A",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"971D",
        x"51E8",
        x"4FFE",
        x"8180",
        x"8191",
        x"81A2",
        x"81B3",
        x"2DE8",
        x"2DF9",
        x"8786",
        x"8797",
        x"8BA0",
        x"8BB1",
        x"CF76",
        x"E011",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"0D8C",
        x"1D9D",
        x"1DAE",
        x"1DBF",
        x"2DE8",
        x"2DF9",
        x"A386",
        x"A397",
        x"A7A0",
        x"A7B1",
        x"CF45",
        x"9628",
        x"E1E0",
        x"940C",
        x"22AC",
        x"2388",
        x"F4A1",
        x"91E0",
        x"00A1",
        x"91F0",
        x"00A2",
        x"9730",
        x"F009",
        x"8210",
        x"1561",
        x"0571",
        x"F019",
        x"2FE6",
        x"2FF7",
        x"8210",
        x"9370",
        x"00A2",
        x"9360",
        x"00A1",
        x"E080",
        x"E090",
        x"9508",
        x"E08B",
        x"E090",
        x"9508",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"972E",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2EA8",
        x"2EB9",
        x"877E",
        x"876D",
        x"2EF4",
        x"2FA8",
        x"2FB9",
        x"921D",
        x"921C",
        x"714E",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"09C5",
        x"9700",
        x"F009",
        x"C118",
        x"2DBF",
        x"71BF",
        x"2E9B",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07C1",
        x"2D2F",
        x"712C",
        x"F409",
        x"C093",
        x"9700",
        x"F099",
        x"3084",
        x"0591",
        x"F009",
        x"C0FE",
        x"EA88",
        x"E093",
        x"940E",
        x"0923",
        x"9700",
        x"F009",
        x"C0F7",
        x"2DE9",
        x"60E8",
        x"2E9E",
        x"9100",
        x"03BA",
        x"9110",
        x"03BB",
        x"C066",
        x"FCF2",
        x"C0E7",
        x"9100",
        x"03BA",
        x"9110",
        x"03BB",
        x"1501",
        x"0511",
        x"F409",
        x"C0E3",
        x"2FA0",
        x"2FB1",
        x"961B",
        x"918C",
        x"971B",
        x"7181",
        x"F009",
        x"C0DB",
        x"FEF3",
        x"C052",
        x"9654",
        x"90CD",
        x"90DC",
        x"9755",
        x"2CE1",
        x"2CF1",
        x"2CEC",
        x"2CFD",
        x"24DD",
        x"24CC",
        x"965A",
        x"918D",
        x"919C",
        x"975B",
        x"E0A0",
        x"E0B0",
        x"2AC8",
        x"2AD9",
        x"2AEA",
        x"2AFB",
        x"2FE0",
        x"2FF1",
        x"8A15",
        x"8A14",
        x"8E13",
        x"8E12",
        x"8E14",
        x"8E15",
        x"8E16",
        x"8E17",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"E021",
        x"2FE8",
        x"2FF9",
        x"8324",
        x"A446",
        x"A457",
        x"A860",
        x"A871",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F0B1",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"940E",
        x"0527",
        x"9700",
        x"F009",
        x"C0A3",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"E081",
        x"1AC8",
        x"08D1",
        x"08E1",
        x"08F1",
        x"86C2",
        x"86D3",
        x"86E4",
        x"86F5",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"012A",
        x"9700",
        x"F009",
        x"C089",
        x"FE93",
        x"C02B",
        x"2FA0",
        x"2FB1",
        x"961B",
        x"921C",
        x"940E",
        x"17F4",
        x"2FE0",
        x"2FF1",
        x"8766",
        x"8777",
        x"8B80",
        x"8B91",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"E081",
        x"8384",
        x"2DF9",
        x"62F0",
        x"2E9F",
        x"C015",
        x"9700",
        x"F009",
        x"C06E",
        x"9100",
        x"03BA",
        x"9110",
        x"03BB",
        x"1501",
        x"0511",
        x"F409",
        x"C062",
        x"2FA0",
        x"2FB1",
        x"961B",
        x"918C",
        x"FD84",
        x"C05C",
        x"FEF1",
        x"C002",
        x"FD80",
        x"C05A",
        x"9120",
        x"03A8",
        x"9130",
        x"03A9",
        x"2FE2",
        x"2FF3",
        x"A546",
        x"A557",
        x"A960",
        x"A971",
        x"2DAA",
        x"2DBB",
        x"965A",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"975D",
        x"9180",
        x"03BA",
        x"9190",
        x"03BB",
        x"965F",
        x"939C",
        x"938E",
        x"975E",
        x"9614",
        x"929C",
        x"2FE0",
        x"2FF1",
        x"8984",
        x"8995",
        x"E0A0",
        x"E0B0",
        x"2FA8",
        x"2FB9",
        x"2799",
        x"2788",
        x"8D42",
        x"8D53",
        x"E060",
        x"E070",
        x"2B84",
        x"2B95",
        x"2BA6",
        x"2BB7",
        x"2DEA",
        x"2DFB",
        x"8786",
        x"8797",
        x"8BA0",
        x"8BB1",
        x"2FE0",
        x"2FF1",
        x"8D84",
        x"8D95",
        x"8DA6",
        x"8DB7",
        x"2DEA",
        x"2DFB",
        x"8782",
        x"8793",
        x"87A4",
        x"87B5",
        x"8216",
        x"8217",
        x"8610",
        x"8611",
        x"EF8F",
        x"8385",
        x"8A16",
        x"8A17",
        x"8E10",
        x"8E11",
        x"8331",
        x"8320",
        x"2FA2",
        x"2FB3",
        x"9616",
        x"918D",
        x"919C",
        x"9717",
        x"8393",
        x"8382",
        x"E080",
        x"C005",
        x"E088",
        x"C003",
        x"E084",
        x"C001",
        x"E087",
        x"E090",
        x"962E",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"9508",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"839C",
        x"838B",
        x"2EA6",
        x"2EB7",
        x"2EE4",
        x"2EF5",
        x"833A",
        x"8329",
        x"2FA2",
        x"2FB3",
        x"921D",
        x"921C",
        x"2FE8",
        x"2FF9",
        x"8162",
        x"8173",
        x"8180",
        x"8191",
        x"940E",
        x"01D8",
        x"9700",
        x"F009",
        x"C18F",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"FD87",
        x"C184",
        x"FF80",
        x"C184",
        x"961A",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"81EB",
        x"81FC",
        x"8146",
        x"8157",
        x"8560",
        x"8571",
        x"1B84",
        x"0B95",
        x"0BA6",
        x"0BB7",
        x"2D4E",
        x"2D5F",
        x"E060",
        x"E070",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F410",
        x"2EE8",
        x"2EF9",
        x"802B",
        x"803C",
        x"E2F0",
        x"0E2F",
        x"1C31",
        x"14E1",
        x"04F1",
        x"F409",
        x"C15C",
        x"81AB",
        x"81BC",
        x"9616",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9719",
        x"2FB7",
        x"2FA6",
        x"2F95",
        x"2F84",
        x"7091",
        x"27AA",
        x"27BB",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F009",
        x"C105",
        x"81EB",
        x"81FC",
        x"8180",
        x"8191",
        x"8135",
        x"2FA8",
        x"2FB9",
        x"9612",
        x"912C",
        x"1732",
        x"F160",
        x"2B45",
        x"2B46",
        x"2B47",
        x"F429",
        x"8566",
        x"8577",
        x"8980",
        x"8991",
        x"C008",
        x"81EB",
        x"81FC",
        x"8942",
        x"8953",
        x"8964",
        x"8975",
        x"940E",
        x"026F",
        x"3062",
        x"0571",
        x"0581",
        x"0591",
        x"F138",
        x"3F6F",
        x"EFBF",
        x"077B",
        x"078B",
        x"079B",
        x"F431",
        x"81EB",
        x"81FC",
        x"8184",
        x"6880",
        x"8384",
        x"C0CD",
        x"81AB",
        x"81BC",
        x"9652",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"9755",
        x"9615",
        x"921C",
        x"81EB",
        x"81FC",
        x"8080",
        x"8091",
        x"8942",
        x"8953",
        x"8964",
        x"8975",
        x"2D88",
        x"2D99",
        x"940E",
        x"059E",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F449",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"6880",
        x"9614",
        x"938C",
        x"C0F9",
        x"81EB",
        x"81FC",
        x"8125",
        x"2E46",
        x"2E57",
        x"2E68",
        x"2E79",
        x"0E42",
        x"1C51",
        x"1C61",
        x"1C71",
        x"2CCE",
        x"2CDF",
        x"2CCD",
        x"24DD",
        x"94C6",
        x"14C1",
        x"04D1",
        x"F409",
        x"C054",
        x"2DA8",
        x"2DB9",
        x"9612",
        x"918C",
        x"E030",
        x"2D4C",
        x"2D5D",
        x"0F42",
        x"1F53",
        x"E090",
        x"1784",
        x"0795",
        x"F420",
        x"2EC8",
        x"2ED9",
        x"1AC2",
        x"0AD3",
        x"2D0C",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D6A",
        x"2D7B",
        x"2DE8",
        x"2DF9",
        x"8181",
        x"940E",
        x"17FF",
        x"81AB",
        x"81BC",
        x"9614",
        x"912C",
        x"9714",
        x"2B89",
        x"F021",
        x"6820",
        x"9614",
        x"932C",
        x"C06D",
        x"FF26",
        x"C01E",
        x"81EB",
        x"81FC",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1984",
        x"0995",
        x"09A6",
        x"09B7",
        x"2D4C",
        x"2D5D",
        x"E060",
        x"E070",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F458",
        x"2F98",
        x"2788",
        x"0F99",
        x"E040",
        x"E052",
        x"2D62",
        x"2D73",
        x"0D8A",
        x"1D9B",
        x"940E",
        x"0099",
        x"81AB",
        x"81BC",
        x"9615",
        x"918C",
        x"9715",
        x"0D8C",
        x"9615",
        x"938C",
        x"2CDC",
        x"24CC",
        x"0CDD",
        x"C073",
        x"81EB",
        x"81FC",
        x"8184",
        x"FF86",
        x"C01A",
        x"8926",
        x"8937",
        x"8D40",
        x"8D51",
        x"E001",
        x"2D62",
        x"2D73",
        x"2DA8",
        x"2DB9",
        x"9611",
        x"918C",
        x"940E",
        x"1809",
        x"81EB",
        x"81FC",
        x"8124",
        x"2B89",
        x"F019",
        x"6820",
        x"8324",
        x"C027",
        x"7B2F",
        x"81AB",
        x"81BC",
        x"9614",
        x"932C",
        x"81EB",
        x"81FC",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1584",
        x"0595",
        x"05A6",
        x"05B7",
        x"F0C9",
        x"9001",
        x"81F0",
        x"2DE0",
        x"E001",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D62",
        x"2D73",
        x"8181",
        x"940E",
        x"17FF",
        x"2B89",
        x"F051",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"6880",
        x"9614",
        x"938C",
        x"E081",
        x"C051",
        x"81EB",
        x"81FC",
        x"8A46",
        x"8A57",
        x"8E60",
        x"8E71",
        x"8185",
        x"5F8F",
        x"8385",
        x"81AB",
        x"81BC",
        x"9616",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9719",
        x"2F84",
        x"2F95",
        x"7091",
        x"E0E0",
        x"E0F2",
        x"1BE8",
        x"0BF9",
        x"2CCE",
        x"2CDF",
        x"15EE",
        x"05FF",
        x"F410",
        x"2ECE",
        x"2EDF",
        x"7051",
        x"2766",
        x"2777",
        x"2F64",
        x"2F75",
        x"5E60",
        x"4F7F",
        x"812B",
        x"813C",
        x"0F62",
        x"1F73",
        x"2D4C",
        x"2D5D",
        x"2D8A",
        x"2D9B",
        x"940E",
        x"0099",
        x"0CAC",
        x"1CBD",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"0D8C",
        x"1D9D",
        x"1DA1",
        x"1DB1",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"81A9",
        x"81BA",
        x"918D",
        x"919C",
        x"9711",
        x"0D8C",
        x"1D9D",
        x"938D",
        x"939C",
        x"18EC",
        x"08FD",
        x"CEA0",
        x"E080",
        x"C003",
        x"E082",
        x"C001",
        x"E087",
        x"E090",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"903F",
        x"902F",
        x"9508",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"839C",
        x"838B",
        x"2EA6",
        x"2EB7",
        x"2EE4",
        x"2EF5",
        x"833A",
        x"8329",
        x"2FA2",
        x"2FB3",
        x"921D",
        x"921C",
        x"2FE8",
        x"2FF9",
        x"8162",
        x"8173",
        x"8180",
        x"8191",
        x"940E",
        x"01D8",
        x"9700",
        x"F009",
        x"C1DD",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"FD87",
        x"C1D2",
        x"FF81",
        x"C1D2",
        x"961A",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"0D4E",
        x"1D5F",
        x"1D61",
        x"1D71",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F410",
        x"2CE1",
        x"2CF1",
        x"802B",
        x"803C",
        x"E2B0",
        x"0E2B",
        x"1C31",
        x"14E1",
        x"04F1",
        x"F409",
        x"C04D",
        x"81EB",
        x"81FC",
        x"8146",
        x"8157",
        x"8560",
        x"8571",
        x"2FB7",
        x"2FA6",
        x"2F95",
        x"2F84",
        x"7091",
        x"27AA",
        x"27BB",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F009",
        x"C153",
        x"9001",
        x"81F0",
        x"2DE0",
        x"81AB",
        x"81BC",
        x"9615",
        x"913C",
        x"9715",
        x"8122",
        x"1732",
        x"F408",
        x"C06A",
        x"2B45",
        x"2B46",
        x"2B47",
        x"F4D1",
        x"961E",
        x"916D",
        x"917D",
        x"918D",
        x"919C",
        x"9751",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F5B9",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F8E",
        x"2F9F",
        x"940E",
        x"043E",
        x"81EB",
        x"81FC",
        x"8766",
        x"8777",
        x"8B80",
        x"8B91",
        x"C00C",
        x"81AB",
        x"81BC",
        x"9652",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9755",
        x"2F8E",
        x"2F9F",
        x"940E",
        x"043E",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F4B9",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"8542",
        x"8553",
        x"8564",
        x"8575",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C14B",
        x"81EB",
        x"81FC",
        x"8782",
        x"8793",
        x"87A4",
        x"87B5",
        x"C144",
        x"81AB",
        x"81BC",
        x"9614",
        x"912C",
        x"9714",
        x"3061",
        x"0571",
        x"0581",
        x"0591",
        x"F429",
        x"2F82",
        x"6880",
        x"9614",
        x"938C",
        x"C13F",
        x"3F6F",
        x"EFBF",
        x"077B",
        x"078B",
        x"079B",
        x"F429",
        x"2F82",
        x"6880",
        x"81EB",
        x"81FC",
        x"C0D6",
        x"81AB",
        x"81BC",
        x"9652",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"9755",
        x"9615",
        x"921C",
        x"81EB",
        x"81FC",
        x"8184",
        x"FF86",
        x"C01C",
        x"8926",
        x"8937",
        x"8D40",
        x"8D51",
        x"9001",
        x"81F0",
        x"2DE0",
        x"E001",
        x"2D62",
        x"2D73",
        x"8181",
        x"940E",
        x"1809",
        x"81AB",
        x"81BC",
        x"9614",
        x"912C",
        x"9714",
        x"2B89",
        x"F021",
        x"6820",
        x"9614",
        x"932C",
        x"C0B0",
        x"7B2F",
        x"81EB",
        x"81FC",
        x"8324",
        x"81AB",
        x"81BC",
        x"908D",
        x"909C",
        x"9711",
        x"9652",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9755",
        x"2D88",
        x"2D99",
        x"940E",
        x"059E",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F431",
        x"81EB",
        x"81FC",
        x"8184",
        x"6880",
        x"8384",
        x"C0EF",
        x"81AB",
        x"81BC",
        x"9615",
        x"912C",
        x"2E46",
        x"2E57",
        x"2E68",
        x"2E79",
        x"0E42",
        x"1C51",
        x"1C61",
        x"1C71",
        x"2CCE",
        x"2CDF",
        x"2CCD",
        x"24DD",
        x"94C6",
        x"14C1",
        x"04D1",
        x"F409",
        x"C051",
        x"2DE8",
        x"2DF9",
        x"8182",
        x"E030",
        x"2D4C",
        x"2D5D",
        x"0F42",
        x"1F53",
        x"E090",
        x"1784",
        x"0795",
        x"F420",
        x"2EC8",
        x"2ED9",
        x"1AC2",
        x"0AD3",
        x"2D0C",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D6A",
        x"2D7B",
        x"2DA8",
        x"2DB9",
        x"9611",
        x"918C",
        x"940E",
        x"1809",
        x"81EB",
        x"81FC",
        x"2B89",
        x"F009",
        x"C058",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1984",
        x"0995",
        x"09A6",
        x"09B7",
        x"2D4C",
        x"2D5D",
        x"E060",
        x"E070",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F4A8",
        x"2F68",
        x"2F79",
        x"2F76",
        x"2766",
        x"0F77",
        x"0D6A",
        x"1D7B",
        x"E040",
        x"E052",
        x"2D82",
        x"2D93",
        x"940E",
        x"0099",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"7B8F",
        x"9614",
        x"938C",
        x"81EB",
        x"81FC",
        x"8185",
        x"0D8C",
        x"8385",
        x"2CDC",
        x"24CC",
        x"0CDD",
        x"C063",
        x"81EB",
        x"81FC",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1584",
        x"0595",
        x"05A6",
        x"05B7",
        x"F119",
        x"8146",
        x"8157",
        x"8560",
        x"8571",
        x"8582",
        x"8593",
        x"85A4",
        x"85B5",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F4B0",
        x"E001",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D62",
        x"2D73",
        x"2DA8",
        x"2DB9",
        x"9611",
        x"918C",
        x"940E",
        x"17FF",
        x"2B89",
        x"F039",
        x"81EB",
        x"81FC",
        x"8184",
        x"6880",
        x"8384",
        x"E081",
        x"C05E",
        x"81AB",
        x"81BC",
        x"9656",
        x"924D",
        x"925D",
        x"926D",
        x"927C",
        x"9759",
        x"9615",
        x"918C",
        x"9715",
        x"5F8F",
        x"9615",
        x"938C",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"2F28",
        x"2F39",
        x"7031",
        x"E040",
        x"E052",
        x"1B42",
        x"0B53",
        x"2CCE",
        x"2CDF",
        x"154E",
        x"055F",
        x"F410",
        x"2EC4",
        x"2ED5",
        x"7091",
        x"27AA",
        x"27BB",
        x"9680",
        x"2D4C",
        x"2D5D",
        x"2D6A",
        x"2D7B",
        x"81AB",
        x"81BC",
        x"0F8A",
        x"1F9B",
        x"940E",
        x"0099",
        x"81EB",
        x"81FC",
        x"8184",
        x"6480",
        x"8384",
        x"0CAC",
        x"1CBD",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"0D8C",
        x"1D9D",
        x"1DA1",
        x"1DB1",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"81A9",
        x"81BA",
        x"918D",
        x"919C",
        x"9711",
        x"0D8C",
        x"1D9D",
        x"938D",
        x"939C",
        x"18EC",
        x"08FD",
        x"CE54",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"6280",
        x"9614",
        x"938C",
        x"E080",
        x"C003",
        x"E082",
        x"C001",
        x"E087",
        x"E090",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"903F",
        x"902F",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"816A",
        x"817B",
        x"8188",
        x"8199",
        x"940E",
        x"01D8",
        x"2F28",
        x"2F39",
        x"9700",
        x"F009",
        x"C054",
        x"818C",
        x"FF85",
        x"C04C",
        x"FF86",
        x"C013",
        x"892E",
        x"893F",
        x"8D48",
        x"8D59",
        x"81E8",
        x"81F9",
        x"E001",
        x"2F6C",
        x"2F7D",
        x"5E60",
        x"4F7F",
        x"8181",
        x"940E",
        x"1809",
        x"2B89",
        x"F5E1",
        x"818C",
        x"7B8F",
        x"838C",
        x"8D4A",
        x"8D5B",
        x"8D6C",
        x"8D7D",
        x"8188",
        x"8199",
        x"940E",
        x"012A",
        x"2F28",
        x"2F39",
        x"9700",
        x"F581",
        x"8D0E",
        x"8D1F",
        x"2FE0",
        x"2FF1",
        x"8583",
        x"6280",
        x"8783",
        x"858A",
        x"859B",
        x"85AC",
        x"85BD",
        x"8F84",
        x"8F95",
        x"8FA6",
        x"8FB7",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8F53",
        x"8F42",
        x"8B75",
        x"8B64",
        x"940E",
        x"17F4",
        x"2FE0",
        x"2FF1",
        x"8B66",
        x"8B77",
        x"8F80",
        x"8F91",
        x"818C",
        x"7D8F",
        x"838C",
        x"81E8",
        x"81F9",
        x"E081",
        x"8384",
        x"8188",
        x"8199",
        x"940E",
        x"01F2",
        x"C007",
        x"E080",
        x"C001",
        x"E081",
        x"E090",
        x"C002",
        x"2F82",
        x"2F93",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"1122",
        x"9700",
        x"F411",
        x"8219",
        x"8218",
        x"91DF",
        x"91CF",
        x"9508",
        x"2388",
        x"F429",
        x"9210",
        x"009E",
        x"E080",
        x"E090",
        x"9508",
        x"E08B",
        x"E090",
        x"9508",
        x"E0AE",
        x"E0B0",
        x"EAEB",
        x"E1F1",
        x"940C",
        x"229C",
        x"879E",
        x"878D",
        x"E040",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"09C5",
        x"9700",
        x"F009",
        x"C045",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07C1",
        x"9700",
        x"F589",
        x"91A0",
        x"03BA",
        x"91B0",
        x"03BB",
        x"9710",
        x"F449",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"8A16",
        x"8A17",
        x"8E10",
        x"8E11",
        x"C027",
        x"961B",
        x"912C",
        x"971B",
        x"FF24",
        x"C020",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"9654",
        x"914D",
        x"915C",
        x"9755",
        x"E060",
        x"E070",
        x"2F64",
        x"2F75",
        x"2755",
        x"2744",
        x"965A",
        x"910D",
        x"911C",
        x"975B",
        x"E020",
        x"E030",
        x"2B40",
        x"2B51",
        x"2B62",
        x"2B73",
        x"8B46",
        x"8B57",
        x"8F60",
        x"8F71",
        x"C005",
        x"3084",
        x"0591",
        x"F411",
        x"E085",
        x"E090",
        x"962E",
        x"E0E4",
        x"940C",
        x"22B8",
        x"E0A4",
        x"E0B0",
        x"E0E7",
        x"E1F2",
        x"940C",
        x"228E",
        x"2E28",
        x"2E39",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"2FA8",
        x"2FB9",
        x"9612",
        x"916D",
        x"917C",
        x"9713",
        x"918D",
        x"919C",
        x"940E",
        x"01D8",
        x"9700",
        x"F009",
        x"C1D7",
        x"2DE2",
        x"2DF3",
        x"8124",
        x"FD27",
        x"C1CE",
        x"8582",
        x"8593",
        x"85A4",
        x"85B5",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F430",
        x"FD21",
        x"C004",
        x"2EC8",
        x"2ED9",
        x"2EEA",
        x"2EFB",
        x"2DA2",
        x"2DB3",
        x"9616",
        x"904D",
        x"905D",
        x"906D",
        x"907C",
        x"9719",
        x"2DE2",
        x"2DF3",
        x"8216",
        x"8217",
        x"8610",
        x"8611",
        x"EF8F",
        x"8385",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F429",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"C139",
        x"8100",
        x"8111",
        x"2FE0",
        x"2FF1",
        x"8082",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"E049",
        x"0C88",
        x"1C99",
        x"1CAA",
        x"1CBB",
        x"954A",
        x"F7D1",
        x"1441",
        x"0451",
        x"0461",
        x"0471",
        x"F409",
        x"C045",
        x"E0F1",
        x"1A4F",
        x"0851",
        x"0861",
        x"0871",
        x"2D9F",
        x"2D8E",
        x"2D7D",
        x"2D6C",
        x"5061",
        x"0971",
        x"0981",
        x"0991",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"940E",
        x"2241",
        x"8329",
        x"833A",
        x"834B",
        x"835C",
        x"2D97",
        x"2D86",
        x"2D75",
        x"2D64",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"940E",
        x"2241",
        x"8169",
        x"817A",
        x"818B",
        x"819C",
        x"1762",
        x"0773",
        x"0784",
        x"0795",
        x"F0D8",
        x"2788",
        x"2799",
        x"27AA",
        x"27BB",
        x"1988",
        x"0999",
        x"09AA",
        x"09BB",
        x"2184",
        x"2195",
        x"21A6",
        x"21B7",
        x"2DE2",
        x"2DF3",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"1AC8",
        x"0AD9",
        x"0AEA",
        x"0AFB",
        x"8942",
        x"8953",
        x"8964",
        x"8975",
        x"C034",
        x"2DA2",
        x"2DB3",
        x"961E",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9751",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F4F9",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"043E",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"3041",
        x"0551",
        x"0561",
        x"0571",
        x"F409",
        x"C0AD",
        x"3F4F",
        x"EFFF",
        x"075F",
        x"076F",
        x"077F",
        x"F409",
        x"C063",
        x"2DE2",
        x"2DF3",
        x"8746",
        x"8757",
        x"8B60",
        x"8B71",
        x"2DA2",
        x"2DB3",
        x"9652",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9755",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F409",
        x"CF67",
        x"C030",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"C08B",
        x"2DA2",
        x"2DB3",
        x"91ED",
        x"91FC",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C07D",
        x"2DA2",
        x"2DB3",
        x"9652",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9755",
        x"9616",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"0D88",
        x"1D99",
        x"1DAA",
        x"1DBB",
        x"2DE2",
        x"2DF3",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"18C8",
        x"08D9",
        x"08EA",
        x"08FB",
        x"148C",
        x"049D",
        x"04AE",
        x"04BF",
        x"F568",
        x"2DE2",
        x"2DF3",
        x"8124",
        x"8180",
        x"8191",
        x"FF21",
        x"C01B",
        x"940E",
        x"043E",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F0B9",
        x"3F4F",
        x"EFFF",
        x"075F",
        x"076F",
        x"077F",
        x"F009",
        x"CFB2",
        x"2DA2",
        x"2DB3",
        x"9614",
        x"918C",
        x"9714",
        x"6880",
        x"9614",
        x"938C",
        x"C098",
        x"940E",
        x"026F",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"CFE9",
        x"2CFB",
        x"2CEA",
        x"2CD9",
        x"2CC8",
        x"2DE2",
        x"2DF3",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"0D8C",
        x"1D9D",
        x"1DAE",
        x"1DBF",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"2C8C",
        x"2C9D",
        x"2CAE",
        x"2CBF",
        x"E039",
        x"94B6",
        x"94A7",
        x"9497",
        x"9487",
        x"953A",
        x"F7D1",
        x"8285",
        x"E0F1",
        x"22DF",
        x"24EE",
        x"24FF",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F409",
        x"CEE0",
        x"2DA2",
        x"2DB3",
        x"918D",
        x"919C",
        x"940E",
        x"059E",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F431",
        x"2DE2",
        x"2DF3",
        x"8184",
        x"6880",
        x"8384",
        x"C079",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"0CC8",
        x"1CD9",
        x"1CEA",
        x"1CFB",
        x"9483",
        x"2DA2",
        x"2DB3",
        x"9615",
        x"928C",
        x"2DE2",
        x"2DF3",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"7091",
        x"27AA",
        x"27BB",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F409",
        x"C047",
        x"8926",
        x"8937",
        x"8D40",
        x"8D51",
        x"16C2",
        x"06D3",
        x"06E4",
        x"06F5",
        x"F1F1",
        x"8184",
        x"2D62",
        x"2D73",
        x"5E60",
        x"4F7F",
        x"2EA6",
        x"2EB7",
        x"FF86",
        x"C016",
        x"9001",
        x"81F0",
        x"2DE0",
        x"E001",
        x"8181",
        x"940E",
        x"1809",
        x"2DA2",
        x"2DB3",
        x"9614",
        x"912C",
        x"9714",
        x"2B89",
        x"F021",
        x"6820",
        x"9614",
        x"932C",
        x"C019",
        x"7B2F",
        x"2DE2",
        x"2DF3",
        x"8324",
        x"2DA2",
        x"2DB3",
        x"91ED",
        x"91FC",
        x"E001",
        x"2D5F",
        x"2D4E",
        x"2D3D",
        x"2D2C",
        x"2D6A",
        x"2D7B",
        x"8181",
        x"940E",
        x"17FF",
        x"2B89",
        x"F039",
        x"2DE2",
        x"2DF3",
        x"8184",
        x"6880",
        x"8384",
        x"E081",
        x"C022",
        x"2DA2",
        x"2DB3",
        x"9656",
        x"92CD",
        x"92DD",
        x"92ED",
        x"92FC",
        x"9759",
        x"2DE2",
        x"2DF3",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"8542",
        x"8553",
        x"8564",
        x"8575",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F450",
        x"8782",
        x"8793",
        x"87A4",
        x"87B5",
        x"8184",
        x"6280",
        x"8384",
        x"C002",
        x"E082",
        x"C001",
        x"E080",
        x"E090",
        x"9624",
        x"E1E2",
        x"940C",
        x"22AA",
        x"E0AE",
        x"E0B0",
        x"EFEB",
        x"E1F3",
        x"940C",
        x"229A",
        x"2EE8",
        x"2EF9",
        x"877E",
        x"876D",
        x"E040",
        x"2F68",
        x"2F79",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"09C5",
        x"9700",
        x"F009",
        x"C048",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2DAE",
        x"2DBF",
        x"9655",
        x"939C",
        x"938E",
        x"9754",
        x"856D",
        x"857E",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"07C1",
        x"9700",
        x"F591",
        x"2DAE",
        x"2DBF",
        x"9652",
        x"91ED",
        x"91FC",
        x"9753",
        x"9730",
        x"F0C9",
        x"8583",
        x"FF84",
        x"C02A",
        x"8944",
        x"8955",
        x"E060",
        x"E070",
        x"2F64",
        x"2F75",
        x"2755",
        x"2744",
        x"8D02",
        x"8D13",
        x"E020",
        x"E030",
        x"2B40",
        x"2B51",
        x"2B62",
        x"2B73",
        x"2DEE",
        x"2DFF",
        x"8346",
        x"8357",
        x"8760",
        x"8771",
        x"2DAE",
        x"2DBF",
        x"91ED",
        x"91FC",
        x"9711",
        x"8186",
        x"8197",
        x"9613",
        x"939C",
        x"938E",
        x"9712",
        x"E060",
        x"E070",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"05E4",
        x"3084",
        x"0591",
        x"F411",
        x"E085",
        x"E090",
        x"962E",
        x"E0E6",
        x"940C",
        x"22B6",
        x"E0AC",
        x"E0B0",
        x"E5EC",
        x"E1F4",
        x"940C",
        x"2298",
        x"2F08",
        x"2F19",
        x"2EC6",
        x"2ED7",
        x"2FE8",
        x"2FF9",
        x"8162",
        x"8173",
        x"8180",
        x"8191",
        x"940E",
        x"01D8",
        x"2EE8",
        x"2EF9",
        x"9700",
        x"F5C9",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2FE0",
        x"2FF1",
        x"8B95",
        x"8B84",
        x"14C1",
        x"04D1",
        x"F439",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"05E4",
        x"C026",
        x"2F80",
        x"2F91",
        x"940E",
        x"0980",
        x"3084",
        x"0591",
        x"F439",
        x"2FE0",
        x"2FF1",
        x"8616",
        x"8617",
        x"8A10",
        x"8A11",
        x"C002",
        x"9700",
        x"F4B1",
        x"2D6C",
        x"2D7D",
        x"2F80",
        x"2F91",
        x"940E",
        x"00A8",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"06AF",
        x"3084",
        x"0591",
        x"F439",
        x"2FE0",
        x"2FF1",
        x"8616",
        x"8617",
        x"8A10",
        x"8A11",
        x"C002",
        x"2EE8",
        x"2EF9",
        x"2D8E",
        x"2D9F",
        x"962C",
        x"E0E8",
        x"940C",
        x"22B4",
        x"E0AE",
        x"E0B0",
        x"EBE1",
        x"E1F4",
        x"940C",
        x"229A",
        x"879E",
        x"878D",
        x"2EE6",
        x"2EF7",
        x"E040",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"09C5",
        x"2F08",
        x"2F19",
        x"9700",
        x"F501",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07C1",
        x"2F08",
        x"2F19",
        x"9700",
        x"F479",
        x"9180",
        x"03BA",
        x"9190",
        x"03BB",
        x"2B89",
        x"F039",
        x"2D6E",
        x"2D7F",
        x"EA88",
        x"E093",
        x"940E",
        x"00A8",
        x"C002",
        x"E006",
        x"E010",
        x"2F80",
        x"2F91",
        x"962E",
        x"E0E6",
        x"940C",
        x"22B6",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"97A4",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"A39C",
        x"A38B",
        x"E041",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"9683",
        x"940E",
        x"09C5",
        x"2F28",
        x"2F39",
        x"9700",
        x"F009",
        x"C08F",
        x"2F8C",
        x"2F9D",
        x"9647",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"A16B",
        x"A17C",
        x"EA88",
        x"E093",
        x"940E",
        x"07C1",
        x"2F28",
        x"2F39",
        x"9700",
        x"F009",
        x"C07D",
        x"91E0",
        x"03BC",
        x"91F0",
        x"03BD",
        x"8583",
        x"FD85",
        x"C074",
        x"91E0",
        x"03BA",
        x"91F0",
        x"03BB",
        x"9730",
        x"F409",
        x"C06A",
        x"8523",
        x"FF20",
        x"C002",
        x"E087",
        x"C066",
        x"88C4",
        x"88D5",
        x"2CE1",
        x"2CF1",
        x"2CEC",
        x"2CFD",
        x"24DD",
        x"24CC",
        x"8D82",
        x"8D93",
        x"E0A0",
        x"E0B0",
        x"2AC8",
        x"2AD9",
        x"2AEA",
        x"2AFB",
        x"FD24",
        x"C009",
        x"EA88",
        x"E093",
        x"940E",
        x"0690",
        x"2F28",
        x"2F39",
        x"9700",
        x"F171",
        x"C04F",
        x"E082",
        x"16C8",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F408",
        x"C041",
        x"E146",
        x"E050",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"0099",
        x"82CF",
        x"86D8",
        x"86E9",
        x"86FA",
        x"E062",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"05E4",
        x"2F28",
        x"2F39",
        x"9700",
        x"F581",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"0980",
        x"2F28",
        x"2F39",
        x"9700",
        x"F409",
        x"CFBA",
        x"3084",
        x"0591",
        x"F259",
        x"C022",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F439",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"01F2",
        x"C018",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"0527",
        x"2F28",
        x"2F39",
        x"9700",
        x"F441",
        x"CFEA",
        x"E082",
        x"C001",
        x"E086",
        x"E090",
        x"C004",
        x"E026",
        x"E030",
        x"2F82",
        x"2F93",
        x"96A4",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"9508",
        x"E1A6",
        x"E0B0",
        x"EAE8",
        x"E1F5",
        x"940C",
        x"228E",
        x"879E",
        x"878D",
        x"E041",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"09C5",
        x"2F28",
        x"2F39",
        x"9700",
        x"F501",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07C1",
        x"2F28",
        x"2F39",
        x"9700",
        x"F069",
        x"3084",
        x"0591",
        x"F461",
        x"91E0",
        x"03BC",
        x"91F0",
        x"03BD",
        x"8583",
        x"FF85",
        x"C008",
        x"E026",
        x"E030",
        x"C002",
        x"E028",
        x"E030",
        x"2F82",
        x"2F93",
        x"C118",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"043E",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F071",
        x"E031",
        x"16C3",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F051",
        x"EF8F",
        x"16C8",
        x"06D8",
        x"06E8",
        x"06F8",
        x"F439",
        x"E081",
        x"C003",
        x"E087",
        x"C001",
        x"E082",
        x"E090",
        x"C0F2",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"012A",
        x"2F28",
        x"2F39",
        x"9700",
        x"F649",
        x"9100",
        x"03A8",
        x"9110",
        x"03A9",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2F80",
        x"2F91",
        x"940E",
        x"059E",
        x"8B6B",
        x"877F",
        x"2F38",
        x"8B9C",
        x"2FA0",
        x"2FB1",
        x"96D2",
        x"910D",
        x"911C",
        x"97D3",
        x"2E20",
        x"2E31",
        x"EFBE",
        x"1A3B",
        x"2FE0",
        x"2FF1",
        x"15E2",
        x"05F3",
        x"F011",
        x"9211",
        x"CFFB",
        x"2F80",
        x"2F91",
        x"960B",
        x"2FE0",
        x"2FF1",
        x"E240",
        x"17E8",
        x"07F9",
        x"F011",
        x"9341",
        x"CFFB",
        x"E22E",
        x"2FE0",
        x"2FF1",
        x"8320",
        x"E180",
        x"8783",
        x"8B2E",
        x"8B3D",
        x"940E",
        x"17F4",
        x"2E46",
        x"2E57",
        x"2E68",
        x"2E79",
        x"2FA0",
        x"2FB1",
        x"9656",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"9759",
        x"965B",
        x"92DC",
        x"92CE",
        x"975A",
        x"2C9F",
        x"2C8E",
        x"24AA",
        x"24BB",
        x"9655",
        x"929C",
        x"928E",
        x"9754",
        x"E240",
        x"E050",
        x"2F60",
        x"2F71",
        x"2F80",
        x"2F91",
        x"9680",
        x"940E",
        x"0099",
        x"892E",
        x"2FE0",
        x"2FF1",
        x"A321",
        x"9180",
        x"03AE",
        x"9190",
        x"03AF",
        x"91A0",
        x"03B0",
        x"91B0",
        x"03B1",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"8140",
        x"893D",
        x"3043",
        x"F469",
        x"A146",
        x"A157",
        x"A560",
        x"A571",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F421",
        x"E080",
        x"E090",
        x"E0A0",
        x"E0B0",
        x"2FE0",
        x"2FF1",
        x"AF93",
        x"AF82",
        x"ABB5",
        x"ABA4",
        x"894B",
        x"855F",
        x"2F63",
        x"897C",
        x"E021",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"8182",
        x"2F94",
        x"893B",
        x"1B93",
        x"1798",
        x"F550",
        x"2FB7",
        x"2FA6",
        x"2F95",
        x"2F84",
        x"9601",
        x"1DA1",
        x"1DB1",
        x"878F",
        x"8B98",
        x"8BA9",
        x"8BBA",
        x"A746",
        x"A757",
        x"AB60",
        x"AB71",
        x"8324",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F8E",
        x"2F9F",
        x"8B2E",
        x"940E",
        x"012A",
        x"2F48",
        x"2F59",
        x"892E",
        x"9700",
        x"F5C1",
        x"2FE0",
        x"2FF1",
        x"15E2",
        x"05F3",
        x"F011",
        x"9211",
        x"CFFB",
        x"854F",
        x"8958",
        x"8969",
        x"897A",
        x"CFCC",
        x"EA88",
        x"E093",
        x"940E",
        x"0923",
        x"2F08",
        x"2F19",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"1501",
        x"0511",
        x"F049",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"940E",
        x"0527",
        x"2F80",
        x"2F91",
        x"C017",
        x"91E0",
        x"03BA",
        x"91F0",
        x"03BB",
        x"E120",
        x"8723",
        x"8A46",
        x"8A57",
        x"8E60",
        x"8E71",
        x"8ED3",
        x"8EC2",
        x"8A95",
        x"8A84",
        x"E021",
        x"2FA8",
        x"2FB9",
        x"9614",
        x"932C",
        x"940E",
        x"01F2",
        x"C001",
        x"2F95",
        x"9666",
        x"E1E2",
        x"940C",
        x"22AA",
        x"E4AF",
        x"E0B0",
        x"EFEB",
        x"E1F6",
        x"940C",
        x"229A",
        x"9660",
        x"AF9F",
        x"AF8E",
        x"9760",
        x"2F06",
        x"2F17",
        x"2F8C",
        x"2F9D",
        x"5B8E",
        x"4F9F",
        x"A79C",
        x"A78B",
        x"E041",
        x"2F6C",
        x"2F7D",
        x"5E69",
        x"4F7F",
        x"2F8C",
        x"2F9D",
        x"5B82",
        x"4F9F",
        x"940E",
        x"09C5",
        x"9700",
        x"F009",
        x"C0DA",
        x"898F",
        x"8D98",
        x"839A",
        x"8389",
        x"9660",
        x"AD6E",
        x"AD7F",
        x"9760",
        x"2F8C",
        x"2F9D",
        x"9647",
        x"940E",
        x"07C1",
        x"9700",
        x"F009",
        x"C0CA",
        x"A5EB",
        x"A5FC",
        x"8583",
        x"FD85",
        x"C0B0",
        x"A589",
        x"A59A",
        x"9700",
        x"F409",
        x"C0A8",
        x"2F68",
        x"2F79",
        x"5F65",
        x"4F7F",
        x"E145",
        x"E050",
        x"2F8C",
        x"2F9D",
        x"968D",
        x"940E",
        x"0099",
        x"E146",
        x"E050",
        x"2F6C",
        x"2F7D",
        x"5E69",
        x"4F7F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"0099",
        x"2F60",
        x"2F71",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"07C1",
        x"2F28",
        x"2F39",
        x"9700",
        x"F409",
        x"C084",
        x"3084",
        x"0591",
        x"F009",
        x"C098",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"0923",
        x"2F28",
        x"2F39",
        x"9700",
        x"F009",
        x"C08E",
        x"88EB",
        x"88FC",
        x"E143",
        x"E050",
        x"2F6C",
        x"2F7D",
        x"5D61",
        x"4F7F",
        x"2D8E",
        x"2D9F",
        x"960D",
        x"940E",
        x"0099",
        x"A58D",
        x"6280",
        x"2DAE",
        x"2DBF",
        x"961B",
        x"938C",
        x"971B",
        x"89EF",
        x"8DF8",
        x"E081",
        x"8384",
        x"961B",
        x"918C",
        x"971B",
        x"FF84",
        x"C061",
        x"8109",
        x"811A",
        x"965A",
        x"914D",
        x"915C",
        x"975B",
        x"9654",
        x"918D",
        x"919C",
        x"9755",
        x"2B48",
        x"2B59",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"059E",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F409",
        x"C053",
        x"2F80",
        x"2F91",
        x"940E",
        x"012A",
        x"2F28",
        x"2F39",
        x"81E9",
        x"81FA",
        x"A902",
        x"A913",
        x"9700",
        x"F009",
        x"C048",
        x"2FA0",
        x"2FB1",
        x"9691",
        x"918C",
        x"328E",
        x"F591",
        x"8120",
        x"818F",
        x"8598",
        x"85A9",
        x"85BA",
        x"3023",
        x"F449",
        x"A146",
        x"A157",
        x"A560",
        x"A571",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F029",
        x"2F58",
        x"2F49",
        x"2F3A",
        x"2F2B",
        x"C004",
        x"E050",
        x"E040",
        x"E030",
        x"E020",
        x"2F85",
        x"2F94",
        x"2FA0",
        x"2FB1",
        x"96DB",
        x"939C",
        x"938E",
        x"97DA",
        x"2F83",
        x"2F92",
        x"96D5",
        x"939C",
        x"938E",
        x"97D4",
        x"E081",
        x"8384",
        x"C008",
        x"E088",
        x"C001",
        x"E084",
        x"E090",
        x"C015",
        x"E086",
        x"E090",
        x"C012",
        x"2F8C",
        x"2F9D",
        x"9647",
        x"940E",
        x"0690",
        x"2F28",
        x"2F39",
        x"9700",
        x"F439",
        x"898F",
        x"8D98",
        x"940E",
        x"01F2",
        x"C004",
        x"E022",
        x"E030",
        x"2F82",
        x"2F93",
        x"5BC1",
        x"4FDF",
        x"E0E6",
        x"940C",
        x"22B6",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"9508",
        x"940E",
        x"1879",
        x"9508",
        x"940E",
        x"1871",
        x"9508",
        x"2F86",
        x"2F97",
        x"2F75",
        x"2F64",
        x"2F53",
        x"2F42",
        x"940E",
        x"1920",
        x"E090",
        x"9508",
        x"2F86",
        x"2F97",
        x"2F75",
        x"2F64",
        x"2F53",
        x"2F42",
        x"940E",
        x"19C4",
        x"E090",
        x"9508",
        x"E080",
        x"E090",
        x"9508",
        x"B387",
        x"6B80",
        x"BB87",
        x"98BE",
        x"9A6C",
        x"B18D",
        x"7F8C",
        x"B98D",
        x"9A6E",
        x"9AC4",
        x"9AC7",
        x"9508",
        x"B98F",
        x"9B77",
        x"CFFE",
        x"B18F",
        x"9508",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD4",
        x"2F15",
        x"2F06",
        x"2EF7",
        x"FF87",
        x"C00A",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E787",
        x"940E",
        x"1827",
        x"3082",
        x"F558",
        x"77CF",
        x"9AC4",
        x"EF8F",
        x"940E",
        x"1822",
        x"98C4",
        x"EF8F",
        x"940E",
        x"1822",
        x"2F8C",
        x"940E",
        x"1822",
        x"2D8F",
        x"940E",
        x"1822",
        x"2F80",
        x"940E",
        x"1822",
        x"2F81",
        x"940E",
        x"1822",
        x"2F8D",
        x"940E",
        x"1822",
        x"34C0",
        x"F021",
        x"34C8",
        x"F021",
        x"E081",
        x"C003",
        x"E985",
        x"C001",
        x"E887",
        x"940E",
        x"1822",
        x"E0CA",
        x"EF8F",
        x"940E",
        x"1822",
        x"FF87",
        x"C002",
        x"50C1",
        x"F7C9",
        x"B7CD",
        x"B7DE",
        x"E0E5",
        x"940C",
        x"22B7",
        x"9AC4",
        x"EF8F",
        x"940E",
        x"1822",
        x"9508",
        x"9180",
        x"03BE",
        x"2388",
        x"F411",
        x"E082",
        x"9508",
        x"E080",
        x"9508",
        x"E0A5",
        x"E0B0",
        x"E7EF",
        x"E1F8",
        x"940C",
        x"229A",
        x"940E",
        x"1816",
        x"E01B",
        x"EF8F",
        x"940E",
        x"1822",
        x"5011",
        x"F7D9",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E480",
        x"940E",
        x"1827",
        x"3081",
        x"F009",
        x"C060",
        x"EA4A",
        x"E051",
        x"E060",
        x"E070",
        x"E488",
        x"940E",
        x"1827",
        x"3081",
        x"F561",
        x"2EEC",
        x"2EFD",
        x"E085",
        x"0EE8",
        x"1CF1",
        x"2F0C",
        x"2F1D",
        x"5F0F",
        x"4F1F",
        x"EF8F",
        x"940E",
        x"1822",
        x"2FE0",
        x"2FF1",
        x"9381",
        x"2F0E",
        x"2F1F",
        x"15EE",
        x"05FF",
        x"F7A9",
        x"818B",
        x"3081",
        x"F009",
        x"C03F",
        x"818C",
        x"3A8A",
        x"F5E1",
        x"EE00",
        x"E21E",
        x"E040",
        x"E050",
        x"E060",
        x"E470",
        x"EE89",
        x"940E",
        x"1827",
        x"2388",
        x"F1D9",
        x"5001",
        x"0911",
        x"1501",
        x"0511",
        x"F791",
        x"C02B",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"EE89",
        x"940E",
        x"1827",
        x"3082",
        x"F420",
        x"E092",
        x"2EF9",
        x"EE99",
        x"C003",
        x"24FF",
        x"94F3",
        x"E491",
        x"EA08",
        x"E611",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F89",
        x"839D",
        x"940E",
        x"1827",
        x"819D",
        x"2388",
        x"F031",
        x"5001",
        x"0911",
        x"1501",
        x"0511",
        x"F781",
        x"C008",
        x"E040",
        x"E052",
        x"E060",
        x"E070",
        x"E580",
        x"940E",
        x"1827",
        x"1181",
        x"2CF1",
        x"92F0",
        x"03BE",
        x"940E",
        x"186C",
        x"E081",
        x"20FF",
        x"F119",
        x"E080",
        x"C021",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E78A",
        x"940E",
        x"1827",
        x"2388",
        x"F769",
        x"2F0C",
        x"2F1D",
        x"5F0F",
        x"4F1F",
        x"EF8F",
        x"940E",
        x"1822",
        x"2FE0",
        x"2FF1",
        x"9381",
        x"2F0E",
        x"2F1F",
        x"15EE",
        x"05FF",
        x"F7A9",
        x"8189",
        x"FF86",
        x"C003",
        x"E02C",
        x"2EF2",
        x"CFD9",
        x"E084",
        x"2EF8",
        x"CFD6",
        x"9625",
        x"E0E6",
        x"940C",
        x"22B6",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F18",
        x"2F09",
        x"9180",
        x"03BE",
        x"FD83",
        x"C007",
        x"E039",
        x"0F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"953A",
        x"F7D1",
        x"E581",
        x"940E",
        x"1827",
        x"2388",
        x"F019",
        x"E0C1",
        x"E0D0",
        x"C023",
        x"E3C0",
        x"E7D5",
        x"EF8F",
        x"940E",
        x"1822",
        x"3F8F",
        x"F421",
        x"9721",
        x"9720",
        x"F7C1",
        x"CFF2",
        x"3F8E",
        x"F781",
        x"2FC1",
        x"2FD0",
        x"E000",
        x"E010",
        x"EF8F",
        x"940E",
        x"1822",
        x"9389",
        x"5F0F",
        x"4F1F",
        x"1501",
        x"E082",
        x"0718",
        x"F7B1",
        x"EF8F",
        x"940E",
        x"1822",
        x"EF8F",
        x"940E",
        x"1822",
        x"E0C0",
        x"E0D0",
        x"940E",
        x"186C",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F18",
        x"2F09",
        x"2EF2",
        x"9180",
        x"03BE",
        x"FD83",
        x"C007",
        x"E0E9",
        x"0F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"95EA",
        x"F7D1",
        x"E581",
        x"940E",
        x"1827",
        x"2388",
        x"F019",
        x"E0C1",
        x"E0D0",
        x"C03B",
        x"E3C0",
        x"E7D5",
        x"EF8F",
        x"940E",
        x"1822",
        x"3F8F",
        x"F421",
        x"9721",
        x"9720",
        x"F7C1",
        x"CFF2",
        x"3F8E",
        x"F781",
        x"20FF",
        x"F429",
        x"2FC1",
        x"2FD0",
        x"E000",
        x"E010",
        x"C009",
        x"E0C0",
        x"E0D1",
        x"EF8F",
        x"940E",
        x"1822",
        x"9721",
        x"9720",
        x"F7D1",
        x"CFF2",
        x"EF8F",
        x"940E",
        x"1822",
        x"9389",
        x"5F0F",
        x"4F1F",
        x"1501",
        x"E081",
        x"0718",
        x"F7B1",
        x"20FF",
        x"F049",
        x"EF8F",
        x"940E",
        x"1822",
        x"EF8F",
        x"940E",
        x"1822",
        x"E0C0",
        x"E0D0",
        x"C009",
        x"E0C0",
        x"E0D1",
        x"EF8F",
        x"940E",
        x"1822",
        x"9721",
        x"9720",
        x"F7D1",
        x"CFEE",
        x"940E",
        x"186C",
        x"2F8C",
        x"2F9D",
        x"B7CD",
        x"B7DE",
        x"E0E5",
        x"940C",
        x"22B7",
        x"E0A2",
        x"E0B0",
        x"ECEA",
        x"E1F9",
        x"940C",
        x"229A",
        x"2F18",
        x"2F09",
        x"9180",
        x"03BE",
        x"FD83",
        x"C007",
        x"E0F9",
        x"0F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"95FA",
        x"F7D1",
        x"E588",
        x"940E",
        x"1827",
        x"2388",
        x"F019",
        x"E081",
        x"E090",
        x"C03F",
        x"EF8F",
        x"940E",
        x"1822",
        x"EF8E",
        x"940E",
        x"1822",
        x"2EE1",
        x"2EF0",
        x"E000",
        x"E010",
        x"2DEE",
        x"2DFF",
        x"9181",
        x"2EEE",
        x"2EFF",
        x"940E",
        x"1822",
        x"5F0F",
        x"4F1F",
        x"1501",
        x"E0F2",
        x"071F",
        x"F799",
        x"E080",
        x"940E",
        x"1822",
        x"E080",
        x"940E",
        x"1822",
        x"EF8F",
        x"940E",
        x"1822",
        x"718F",
        x"3085",
        x"F6D1",
        x"EE08",
        x"EF1D",
        x"EF8F",
        x"940E",
        x"1822",
        x"3F8F",
        x"F049",
        x"1501",
        x"0511",
        x"F019",
        x"5001",
        x"0911",
        x"CFF5",
        x"E081",
        x"E090",
        x"C006",
        x"E081",
        x"E090",
        x"1501",
        x"0511",
        x"F009",
        x"E080",
        x"8389",
        x"839A",
        x"940E",
        x"186C",
        x"819A",
        x"8189",
        x"9622",
        x"E0E6",
        x"940C",
        x"22B6",
        x"93CF",
        x"93DF",
        x"9AC3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"B389",
        x"9380",
        x"00A3",
        x"9AC0",
        x"9180",
        x"00A3",
        x"2F98",
        x"7190",
        x"FD84",
        x"C002",
        x"9380",
        x"00A4",
        x"9180",
        x"00A4",
        x"7087",
        x"3081",
        x"F409",
        x"C14E",
        x"F038",
        x"3082",
        x"F409",
        x"C11C",
        x"3083",
        x"F409",
        x"C12C",
        x"C1A3",
        x"2399",
        x"F009",
        x"C1A0",
        x"98C3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"B389",
        x"9380",
        x"00A5",
        x"9AC0",
        x"9120",
        x"00A5",
        x"2F82",
        x"7988",
        x"3180",
        x"F451",
        x"2F82",
        x"9582",
        x"9586",
        x"7087",
        x"E090",
        x"9390",
        x"0064",
        x"9380",
        x"0063",
        x"792F",
        x"2F82",
        x"7F80",
        x"3280",
        x"F459",
        x"2F82",
        x"9586",
        x"9586",
        x"7083",
        x"E090",
        x"9390",
        x"0064",
        x"9380",
        x"0063",
        x"7F23",
        x"C006",
        x"2322",
        x"F409",
        x"C132",
        x"3021",
        x"F409",
        x"C149",
        x"3022",
        x"F409",
        x"C149",
        x"3024",
        x"F409",
        x"C149",
        x"3025",
        x"F409",
        x"C149",
        x"3028",
        x"F409",
        x"C149",
        x"3120",
        x"F409",
        x"C149",
        x"3121",
        x"F409",
        x"C149",
        x"3122",
        x"F409",
        x"C149",
        x"3123",
        x"F409",
        x"C149",
        x"3127",
        x"F409",
        x"C149",
        x"3124",
        x"F409",
        x"C149",
        x"3125",
        x"F409",
        x"C149",
        x"3126",
        x"F409",
        x"C149",
        x"3220",
        x"F481",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"02A8",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"E081",
        x"9380",
        x"03FF",
        x"E082",
        x"9380",
        x"00A4",
        x"C039",
        x"3221",
        x"F429",
        x"9210",
        x"03FF",
        x"9210",
        x"03FA",
        x"C032",
        x"3222",
        x"F451",
        x"9180",
        x"03BF",
        x"E090",
        x"9390",
        x"046F",
        x"9380",
        x"046E",
        x"E2C1",
        x"E1DE",
        x"C0FA",
        x"3223",
        x"F451",
        x"9180",
        x"03BF",
        x"E090",
        x"9390",
        x"046F",
        x"9380",
        x"046E",
        x"E6CC",
        x"E1DE",
        x"C0EE",
        x"332F",
        x"F409",
        x"C118",
        x"3420",
        x"F4C1",
        x"9180",
        x"02A8",
        x"7083",
        x"9380",
        x"03F9",
        x"9180",
        x"02A9",
        x"9190",
        x"02AA",
        x"91A0",
        x"02AB",
        x"91B0",
        x"02AC",
        x"9380",
        x"03FB",
        x"9390",
        x"03FC",
        x"93A0",
        x"03FD",
        x"93B0",
        x"03FE",
        x"E0C0",
        x"E0D0",
        x"C0D1",
        x"3421",
        x"F489",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"03BF",
        x"7083",
        x"E090",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"5480",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8585",
        x"C0A5",
        x"E0C0",
        x"E0D0",
        x"3422",
        x"F409",
        x"C0A8",
        x"3423",
        x"F409",
        x"C0A8",
        x"3424",
        x"F409",
        x"C0A8",
        x"3425",
        x"F409",
        x"C0A8",
        x"3426",
        x"F409",
        x"C0A8",
        x"3427",
        x"F409",
        x"C0A8",
        x"3820",
        x"F449",
        x"E080",
        x"940E",
        x"17F9",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"03BE",
        x"C02D",
        x"3E20",
        x"F429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E28C",
        x"C026",
        x"3E21",
        x"F431",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"02A6",
        x"C01E",
        x"3F20",
        x"F431",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"02A7",
        x"C016",
        x"3F21",
        x"F469",
        x"9160",
        x"03BF",
        x"9360",
        x"02A7",
        x"EF8F",
        x"E090",
        x"940E",
        x"2350",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"C007",
        x"3F2D",
        x"F451",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"00A4",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"C06D",
        x"3F2E",
        x"F009",
        x"C06A",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0060",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9180",
        x"0060",
        x"9580",
        x"9380",
        x"0060",
        x"C05B",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"91E0",
        x"03FF",
        x"E0F0",
        x"55E8",
        x"4FFD",
        x"8180",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9180",
        x"03FF",
        x"5F8F",
        x"9380",
        x"03FF",
        x"C078",
        x"2399",
        x"F009",
        x"C075",
        x"98C3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"B389",
        x"9380",
        x"00A5",
        x"9AC0",
        x"9180",
        x"03FF",
        x"2FE8",
        x"E0F0",
        x"55E8",
        x"4FFD",
        x"9190",
        x"00A5",
        x"8390",
        x"5F8F",
        x"9380",
        x"03FF",
        x"E081",
        x"9380",
        x"03FA",
        x"C05D",
        x"2399",
        x"F009",
        x"C05A",
        x"98C3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"B389",
        x"9380",
        x"00A5",
        x"9AC0",
        x"9180",
        x"00A5",
        x"9380",
        x"03BF",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"03BF",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"C044",
        x"EACF",
        x"E1DC",
        x"C011",
        x"E1C8",
        x"E2D1",
        x"C00E",
        x"ECC8",
        x"E1DF",
        x"C00B",
        x"E1C7",
        x"E2D0",
        x"C008",
        x"EDCE",
        x"E2D0",
        x"C005",
        x"E7CB",
        x"E2D0",
        x"C002",
        x"EEC9",
        x"E2D0",
        x"9720",
        x"F171",
        x"2FEC",
        x"2FFD",
        x"9509",
        x"C02A",
        x"ECCA",
        x"E1DC",
        x"CFF7",
        x"E3CD",
        x"E1DD",
        x"CFF4",
        x"E4CA",
        x"E1DD",
        x"CFF1",
        x"E5C7",
        x"E1DD",
        x"CFEE",
        x"E6C4",
        x"E1DD",
        x"CFEB",
        x"EAC0",
        x"E1DE",
        x"CFE8",
        x"E7C8",
        x"E1DD",
        x"CFE5",
        x"E7CA",
        x"E1DF",
        x"CFE2",
        x"E9C7",
        x"E1DD",
        x"CFDF",
        x"EAC3",
        x"E1DD",
        x"CFDC",
        x"EBC5",
        x"E1DE",
        x"CFD9",
        x"EACF",
        x"E1DD",
        x"CFD6",
        x"ECC2",
        x"E1DE",
        x"CFD3",
        x"E5C1",
        x"E2D1",
        x"CFD0",
        x"91DF",
        x"91CF",
        x"9508",
        x"2F48",
        x"9120",
        x"0063",
        x"9130",
        x"0064",
        x"2B23",
        x"F439",
        x"EA68",
        x"E072",
        x"E780",
        x"E094",
        x"940E",
        x"0BD9",
        x"C03D",
        x"9210",
        x"0064",
        x"9210",
        x"0063",
        x"9120",
        x"0690",
        x"9130",
        x"0691",
        x"2B23",
        x"F419",
        x"E021",
        x"E030",
        x"C011",
        x"9120",
        x"08B0",
        x"9130",
        x"08B1",
        x"2B23",
        x"F419",
        x"E022",
        x"E030",
        x"C008",
        x"9120",
        x"0AD0",
        x"9130",
        x"0AD1",
        x"2B23",
        x"F431",
        x"E023",
        x"E030",
        x"9330",
        x"0064",
        x"9320",
        x"0063",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"1618",
        x"0619",
        x"F494",
        x"E260",
        x"E072",
        x"940E",
        x"2230",
        x"EA68",
        x"E072",
        x"5980",
        x"4F9B",
        x"940E",
        x"0BD9",
        x"9700",
        x"F441",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"6280",
        x"C002",
        x"E182",
        x"E090",
        x"6480",
        x"9508",
        x"9210",
        x"03F8",
        x"EA86",
        x"E090",
        x"9390",
        x"0D35",
        x"9380",
        x"0D34",
        x"E348",
        x"E050",
        x"EF6F",
        x"E070",
        x"EC80",
        x"E093",
        x"940E",
        x"2326",
        x"E080",
        x"940E",
        x"119B",
        x"E062",
        x"E07D",
        x"E080",
        x"940E",
        x"0BC0",
        x"9210",
        x"0471",
        x"9210",
        x"0470",
        x"9210",
        x"0691",
        x"9210",
        x"0690",
        x"9210",
        x"08B1",
        x"9210",
        x"08B0",
        x"9210",
        x"0AD1",
        x"9210",
        x"0AD0",
        x"9508",
        x"EAE8",
        x"E0F2",
        x"9001",
        x"2000",
        x"F7E9",
        x"9731",
        x"5AE8",
        x"40F2",
        x"EAA8",
        x"E0B2",
        x"EF6F",
        x"EF7F",
        x"EF2F",
        x"EF3F",
        x"E080",
        x"E090",
        x"178E",
        x"079F",
        x"F139",
        x"3F2F",
        x"EF4F",
        x"0734",
        x"F489",
        x"914D",
        x"334F",
        x"F039",
        x"324A",
        x"F029",
        x"354C",
        x"F031",
        x"324F",
        x"F431",
        x"C003",
        x"2F28",
        x"2F39",
        x"C002",
        x"2F68",
        x"2F79",
        x"9601",
        x"CFE8",
        x"3F6F",
        x"EF8F",
        x"0778",
        x"F0D1",
        x"2FE6",
        x"2FF7",
        x"55E8",
        x"4FFD",
        x"8210",
        x"5567",
        x"4F7D",
        x"E140",
        x"E050",
        x"EF81",
        x"E09C",
        x"940E",
        x"2337",
        x"9508",
        x"3F2F",
        x"4F3F",
        x"F759",
        x"E140",
        x"E050",
        x"E768",
        x"E070",
        x"EF81",
        x"E09C",
        x"940E",
        x"2305",
        x"9508",
        x"E140",
        x"E050",
        x"EA68",
        x"E072",
        x"EF81",
        x"E09C",
        x"940E",
        x"2337",
        x"9210",
        x"02A8",
        x"9508",
        x"940E",
        x"1C5E",
        x"EA68",
        x"E072",
        x"E588",
        x"E094",
        x"940E",
        x"13F5",
        x"9380",
        x"0CF0",
        x"98C3",
        x"2388",
        x"F031",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0CF0",
        x"6480",
        x"C003",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"E060",
        x"E074",
        x"E588",
        x"E094",
        x"940E",
        x"1456",
        x"9380",
        x"0CF0",
        x"2388",
        x"F421",
        x"9180",
        x"0409",
        x"2388",
        x"F439",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0CF0",
        x"6480",
        x"C050",
        x"E069",
        x"E074",
        x"EF81",
        x"E09C",
        x"940E",
        x"21BF",
        x"2B89",
        x"F319",
        x"E0C9",
        x"E0D4",
        x"9009",
        x"2000",
        x"F7E9",
        x"50CA",
        x"40D4",
        x"2F0C",
        x"9110",
        x"0408",
        x"2F81",
        x"7180",
        x"2EF8",
        x"FF14",
        x"C005",
        x"E38C",
        x"9380",
        x"02A8",
        x"E081",
        x"C001",
        x"E080",
        x"2799",
        x"FD87",
        x"9590",
        x"E069",
        x"E074",
        x"5588",
        x"4F9D",
        x"940E",
        x"232E",
        x"20FF",
        x"F059",
        x"2FEC",
        x"27FF",
        x"FDE7",
        x"95F0",
        x"55E8",
        x"4FFD",
        x"E38E",
        x"8381",
        x"8212",
        x"2F0C",
        x"5F0E",
        x"2F80",
        x"2799",
        x"FD87",
        x"9590",
        x"2FE8",
        x"2FF9",
        x"55E8",
        x"4FFD",
        x"8311",
        x"2FE8",
        x"2FF9",
        x"55E6",
        x"4FFD",
        x"9180",
        x"0400",
        x"9190",
        x"0401",
        x"91A0",
        x"0402",
        x"91B0",
        x"0403",
        x"8380",
        x"8391",
        x"83A2",
        x"83B3",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"B7CD",
        x"B7DE",
        x"E0E5",
        x"940C",
        x"22B7",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"11A5",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"15A2",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"14E7",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"EAE8",
        x"E0F2",
        x"9001",
        x"2000",
        x"F7E9",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"2F6E",
        x"2F7F",
        x"EA88",
        x"E092",
        x"940E",
        x"16F5",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"E081",
        x"940E",
        x"1BE8",
        x"9380",
        x"0CF0",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"3084",
        x"0591",
        x"F444",
        x"E166",
        x"E070",
        x"940E",
        x"2230",
        x"5080",
        x"4F9C",
        x"940E",
        x"09BE",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0CF0",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E086",
        x"940E",
        x"1BE8",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E182",
        x"940E",
        x"1BE8",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"EBE5",
        x"E1FD",
        x"940C",
        x"2294",
        x"9100",
        x"0063",
        x"9110",
        x"0064",
        x"2F80",
        x"2F91",
        x"E260",
        x"E072",
        x"940E",
        x"2230",
        x"2FC8",
        x"2FD9",
        x"59C0",
        x"4FDB",
        x"853A",
        x"852B",
        x"859C",
        x"858D",
        x"9330",
        x"02A8",
        x"9320",
        x"02A9",
        x"9390",
        x"02AA",
        x"9380",
        x"02AB",
        x"9160",
        x"0D04",
        x"E070",
        x"E080",
        x"E090",
        x"852E",
        x"853F",
        x"8948",
        x"8959",
        x"5022",
        x"0931",
        x"0941",
        x"0951",
        x"940E",
        x"226A",
        x"2E82",
        x"2E93",
        x"2EA4",
        x"2EB5",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"9180",
        x"0D2C",
        x"9190",
        x"0D2D",
        x"91A0",
        x"0D2E",
        x"91B0",
        x"0D2F",
        x"0D88",
        x"1D99",
        x"1DAA",
        x"1DBB",
        x"9380",
        x"02AC",
        x"9390",
        x"02AD",
        x"93A0",
        x"02AE",
        x"93B0",
        x"02AF",
        x"813E",
        x"812F",
        x"8598",
        x"8589",
        x"9330",
        x"02B0",
        x"9320",
        x"02B1",
        x"9390",
        x"02B2",
        x"9380",
        x"02B3",
        x"2F80",
        x"2F91",
        x"E166",
        x"E070",
        x"940E",
        x"2230",
        x"5080",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8580",
        x"738F",
        x"9380",
        x"02B4",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"22B0",
        x"E0A2",
        x"E0B0",
        x"E2E7",
        x"E1FE",
        x"940C",
        x"229E",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"2230",
        x"5980",
        x"4F9B",
        x"9120",
        x"046E",
        x"9130",
        x"046F",
        x"2B23",
        x"F431",
        x"E020",
        x"E031",
        x"9330",
        x"046F",
        x"9320",
        x"046E",
        x"9140",
        x"046E",
        x"9150",
        x"046F",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"EA68",
        x"E072",
        x"940E",
        x"0D32",
        x"9120",
        x"0063",
        x"9130",
        x"0064",
        x"1612",
        x"0613",
        x"F484",
        x"9700",
        x"F471",
        x"9140",
        x"046E",
        x"9150",
        x"046F",
        x"8129",
        x"813A",
        x"1742",
        x"0753",
        x"F029",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E680",
        x"C004",
        x"98C3",
        x"EF9F",
        x"BB9A",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"22BA",
        x"E0A2",
        x"E0B0",
        x"E7E2",
        x"E1FE",
        x"940C",
        x"229E",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"2230",
        x"5980",
        x"4F9B",
        x"9120",
        x"046E",
        x"9130",
        x"046F",
        x"2B23",
        x"F431",
        x"E020",
        x"E031",
        x"9330",
        x"046F",
        x"9320",
        x"046E",
        x"98C3",
        x"EF2F",
        x"BB2A",
        x"9140",
        x"046E",
        x"9150",
        x"046F",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"EA68",
        x"E072",
        x"940E",
        x"0F03",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"22BA",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"2230",
        x"98C3",
        x"EF2F",
        x"BB2A",
        x"5980",
        x"4F9B",
        x"940E",
        x"118E",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"14E7",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"2230",
        x"9140",
        x"02A8",
        x"9150",
        x"02A9",
        x"9160",
        x"02AA",
        x"9170",
        x"02AB",
        x"98C3",
        x"EF2F",
        x"BB2A",
        x"5980",
        x"4F9B",
        x"940E",
        x"1201",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"9180",
        x"0061",
        x"9190",
        x"0062",
        x"17C8",
        x"07D9",
        x"F419",
        x"E080",
        x"E090",
        x"C023",
        x"FD97",
        x"C004",
        x"ED80",
        x"E09A",
        x"940E",
        x"118E",
        x"EF8F",
        x"EF9F",
        x"9390",
        x"0062",
        x"9380",
        x"0061",
        x"FDD7",
        x"CFEF",
        x"2F8C",
        x"2F9D",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"2F68",
        x"2F79",
        x"5460",
        x"4F7C",
        x"E043",
        x"ED80",
        x"E09A",
        x"940E",
        x"0BD9",
        x"9700",
        x"F421",
        x"93D0",
        x"0062",
        x"93C0",
        x"0061",
        x"91DF",
        x"91CF",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"1EDF",
        x"9380",
        x"0CF0",
        x"2388",
        x"F011",
        x"6480",
        x"C029",
        x"2F8C",
        x"2F9D",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"2F08",
        x"2F19",
        x"5400",
        x"4F1C",
        x"ECC0",
        x"E0D3",
        x"170C",
        x"071D",
        x"F051",
        x"E04E",
        x"E050",
        x"2F6C",
        x"2F7D",
        x"2F80",
        x"2F91",
        x"940E",
        x"2317",
        x"2B89",
        x"F079",
        x"962E",
        x"E083",
        x"3FC8",
        x"07D8",
        x"F771",
        x"E080",
        x"E094",
        x"940E",
        x"09BE",
        x"9180",
        x"0408",
        x"2FE0",
        x"2FF1",
        x"8785",
        x"C001",
        x"E48A",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"E5E5",
        x"E1FF",
        x"940C",
        x"229E",
        x"E66C",
        x"E070",
        x"EA88",
        x"E092",
        x"940E",
        x"22FB",
        x"E142",
        x"EA68",
        x"E072",
        x"E780",
        x"E094",
        x"940E",
        x"0BD9",
        x"9380",
        x"0CF0",
        x"2388",
        x"F481",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E348",
        x"E050",
        x"EC60",
        x"E073",
        x"E780",
        x"E094",
        x"940E",
        x"0F03",
        x"E780",
        x"E094",
        x"940E",
        x"118E",
        x"9622",
        x"E0E2",
        x"940C",
        x"22BA",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"9100",
        x"02A8",
        x"7003",
        x"E010",
        x"2F80",
        x"2F91",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"2FC8",
        x"2FD9",
        x"54C0",
        x"4FDC",
        x"E08E",
        x"2FEC",
        x"2FFD",
        x"9211",
        x"958A",
        x"F7E9",
        x"E04D",
        x"E050",
        x"EA69",
        x"E072",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"2337",
        x"2F80",
        x"2F91",
        x"940E",
        x"1F13",
        x"2F18",
        x"3480",
        x"F040",
        x"E04E",
        x"E050",
        x"EF6F",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"2326",
        x"940E",
        x"1F4F",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"BB1B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"9140",
        x"03FB",
        x"9150",
        x"03FC",
        x"9160",
        x"03FD",
        x"9170",
        x"03FE",
        x"2F76",
        x"2F65",
        x"2F54",
        x"2744",
        x"ED80",
        x"E09A",
        x"940E",
        x"1201",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"ECEE",
        x"E1FF",
        x"940C",
        x"229E",
        x"9120",
        x"03F9",
        x"E030",
        x"2F82",
        x"2F93",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"5480",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8585",
        x"3F8F",
        x"F169",
        x"2F82",
        x"2F93",
        x"940E",
        x"1EDF",
        x"940E",
        x"1FB7",
        x"2388",
        x"F4A9",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E040",
        x"E051",
        x"EA68",
        x"E072",
        x"ED80",
        x"E09A",
        x"940E",
        x"0D32",
        x"2F28",
        x"2388",
        x"F439",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"C015",
        x"E429",
        x"9180",
        x"03F9",
        x"E090",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"2FE8",
        x"2FF9",
        x"54E0",
        x"4FFC",
        x"EF8F",
        x"8785",
        x"6420",
        x"C001",
        x"E429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"BB2B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"22BA",
        x"E0A2",
        x"E0B0",
        x"E1ED",
        x"E2F0",
        x"940C",
        x"229E",
        x"9120",
        x"03F9",
        x"E030",
        x"2F82",
        x"2F93",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"5480",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8585",
        x"3F8F",
        x"F409",
        x"C041",
        x"FF80",
        x"C005",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E48A",
        x"C022",
        x"2F82",
        x"2F93",
        x"940E",
        x"1EDF",
        x"940E",
        x"1FB7",
        x"2388",
        x"F4E1",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E040",
        x"E051",
        x"EA68",
        x"E072",
        x"ED80",
        x"E09A",
        x"940E",
        x"0F03",
        x"2F28",
        x"2388",
        x"F471",
        x"ED80",
        x"E09A",
        x"940E",
        x"1122",
        x"2F28",
        x"2388",
        x"F439",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"C01B",
        x"E429",
        x"9180",
        x"03F9",
        x"E090",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"2FE8",
        x"2FF9",
        x"54E0",
        x"4FFC",
        x"EF8F",
        x"8785",
        x"98C3",
        x"BB8A",
        x"E480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"C001",
        x"E429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"BB2B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"22BA",
        x"E0A2",
        x"E0B0",
        x"E8E1",
        x"E2F0",
        x"940C",
        x"229A",
        x"E660",
        x"E070",
        x"EA88",
        x"E092",
        x"940E",
        x"22FB",
        x"E041",
        x"EA68",
        x"E072",
        x"E780",
        x"E094",
        x"940E",
        x"0BD9",
        x"9380",
        x"0CF0",
        x"2388",
        x"F499",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E348",
        x"E050",
        x"EC60",
        x"E073",
        x"E780",
        x"E094",
        x"940E",
        x"0D32",
        x"9380",
        x"0CF0",
        x"E780",
        x"E094",
        x"940E",
        x"118E",
        x"C008",
        x"E348",
        x"E050",
        x"EF6F",
        x"E070",
        x"EC80",
        x"E093",
        x"940E",
        x"2326",
        x"EC9D",
        x"2EE9",
        x"E093",
        x"2EF9",
        x"E000",
        x"E010",
        x"2DEE",
        x"2DFF",
        x"8180",
        x"3F8F",
        x"F451",
        x"E04E",
        x"E050",
        x"EF6F",
        x"E070",
        x"2D8E",
        x"2D9F",
        x"970D",
        x"940E",
        x"2326",
        x"C006",
        x"2F80",
        x"2F91",
        x"940E",
        x"1F13",
        x"FD86",
        x"CFF0",
        x"5F0F",
        x"4F1F",
        x"E0FE",
        x"0EEF",
        x"1CF1",
        x"3004",
        x"0511",
        x"F719",
        x"940E",
        x"1F4F",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E6",
        x"940C",
        x"22B6",
        x"940E",
        x"1F4F",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"93CF",
        x"93DF",
        x"91C0",
        x"03BF",
        x"70C3",
        x"E0D0",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1EDF",
        x"ED80",
        x"E09A",
        x"940E",
        x"118E",
        x"EF8F",
        x"EF9F",
        x"9390",
        x"0062",
        x"9380",
        x"0061",
        x"2F8C",
        x"2F9D",
        x"E06E",
        x"E070",
        x"940E",
        x"2230",
        x"E04E",
        x"E050",
        x"EF6F",
        x"E070",
        x"5480",
        x"4F9C",
        x"940E",
        x"2326",
        x"940E",
        x"1F4F",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"91DF",
        x"91CF",
        x"9508",
        x"93CF",
        x"93DF",
        x"ECED",
        x"E0F3",
        x"E050",
        x"8180",
        x"3F8F",
        x"F0C9",
        x"E080",
        x"E090",
        x"2F2E",
        x"2F3F",
        x"502D",
        x"0931",
        x"2F45",
        x"0F48",
        x"2FC2",
        x"2FD3",
        x"0FC8",
        x"1FD9",
        x"8168",
        x"2366",
        x"F059",
        x"9601",
        x"308D",
        x"0591",
        x"F039",
        x"2FA4",
        x"E0B0",
        x"55A8",
        x"4FBD",
        x"936C",
        x"CFED",
        x"2F45",
        x"2FA4",
        x"E0B0",
        x"55A8",
        x"4FBD",
        x"921C",
        x"E051",
        x"0F54",
        x"963E",
        x"E084",
        x"30E5",
        x"07F8",
        x"F6B9",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"91DF",
        x"91CF",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E5E7",
        x"E2F1",
        x"940C",
        x"2298",
        x"9180",
        x"046E",
        x"9190",
        x"046F",
        x"2B89",
        x"F449",
        x"9180",
        x"03FA",
        x"2388",
        x"F429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E488",
        x"C050",
        x"9180",
        x"02A8",
        x"9190",
        x"02A9",
        x"3485",
        x"E522",
        x"0792",
        x"F0C1",
        x"3485",
        x"4597",
        x"F009",
        x"C048",
        x"9180",
        x"02AA",
        x"E090",
        x"9120",
        x"02AB",
        x"2EE8",
        x"2EF9",
        x"0EE2",
        x"1CF1",
        x"EA0C",
        x"E012",
        x"EAC8",
        x"E0D2",
        x"2F28",
        x"2F39",
        x"5A28",
        x"4032",
        x"2EC2",
        x"2ED3",
        x"C01C",
        x"9180",
        x"02AA",
        x"E090",
        x"9120",
        x"02AB",
        x"2F08",
        x"2F19",
        x"0F02",
        x"1D11",
        x"EAC8",
        x"E0D2",
        x"2FE8",
        x"2FF9",
        x"5AE8",
        x"40F2",
        x"2EEE",
        x"2EFF",
        x"2D8E",
        x"2D9F",
        x"0F8C",
        x"1F9D",
        x"1780",
        x"0791",
        x"F4A0",
        x"940E",
        x"2348",
        x"9389",
        x"CFF5",
        x"2D8C",
        x"2D9D",
        x"0F8C",
        x"1F9D",
        x"158E",
        x"059F",
        x"F448",
        x"2FE0",
        x"2FF1",
        x"9161",
        x"2F0E",
        x"2F1F",
        x"940E",
        x"2350",
        x"9621",
        x"CFF0",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"B7CD",
        x"B7DE",
        x"E0E8",
        x"940C",
        x"22B4",
        x"93CF",
        x"93DF",
        x"2FA6",
        x"2FB7",
        x"2FE8",
        x"2FF9",
        x"2FC6",
        x"2FD7",
        x"9139",
        x"2F6C",
        x"2F7D",
        x"2333",
        x"F429",
        x"E040",
        x"E050",
        x"E020",
        x"E030",
        x"C01E",
        x"2FC8",
        x"2FD9",
        x"9129",
        x"2F8C",
        x"2F9D",
        x"322A",
        x"F3A1",
        x"1723",
        x"F339",
        x"332F",
        x"F329",
        x"E080",
        x"C02F",
        x"8180",
        x"328A",
        x"F491",
        x"2F8E",
        x"2F9F",
        x"9601",
        x"8121",
        x"2322",
        x"F129",
        x"2F2A",
        x"2F3B",
        x"5F2F",
        x"4F3F",
        x"2F48",
        x"2F59",
        x"2FE8",
        x"2FF9",
        x"919C",
        x"2399",
        x"F761",
        x"C010",
        x"1789",
        x"F011",
        x"338F",
        x"F429",
        x"2F8E",
        x"2F9F",
        x"9601",
        x"9611",
        x"CFF1",
        x"2FA2",
        x"2FB3",
        x"5F2F",
        x"4F3F",
        x"2F84",
        x"2F95",
        x"CFEA",
        x"9121",
        x"322A",
        x"F3E9",
        x"E081",
        x"E090",
        x"2322",
        x"F021",
        x"E080",
        x"C002",
        x"E081",
        x"E090",
        x"91DF",
        x"91CF",
        x"9508",
        x"E020",
        x"EE31",
        x"E040",
        x"E050",
        x"E060",
        x"EE71",
        x"E080",
        x"E090",
        x"940E",
        x"0095",
        x"940E",
        x"0064",
        x"EF8F",
        x"9380",
        x"02A7",
        x"940E",
        x"1816",
        x"940E",
        x"1C35",
        x"9478",
        x"E180",
        x"BF89",
        x"B608",
        x"FE04",
        x"CFFD",
        x"B788",
        x"6180",
        x"BF88",
        x"940E",
        x"1A22",
        x"CFF7",
        x"2400",
        x"2755",
        x"C004",
        x"0E08",
        x"1F59",
        x"0F88",
        x"1F99",
        x"9700",
        x"F029",
        x"9576",
        x"9567",
        x"F3B8",
        x"0571",
        x"F7B9",
        x"2D80",
        x"2F95",
        x"9508",
        x"E2A1",
        x"2E1A",
        x"1BAA",
        x"1BBB",
        x"2FEA",
        x"2FFB",
        x"C00D",
        x"1FAA",
        x"1FBB",
        x"1FEE",
        x"1FFF",
        x"17A2",
        x"07B3",
        x"07E4",
        x"07F5",
        x"F020",
        x"1BA2",
        x"0BB3",
        x"0BE4",
        x"0BF5",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"941A",
        x"F769",
        x"9560",
        x"9570",
        x"9580",
        x"9590",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"9468",
        x"1000",
        x"94E8",
        x"E0A0",
        x"E0B0",
        x"E7E1",
        x"E2F2",
        x"940C",
        x"2296",
        x"EFEF",
        x"F9E7",
        x"2EA2",
        x"2EB3",
        x"2EC4",
        x"2ED5",
        x"235E",
        x"0F55",
        x"08EE",
        x"2CFE",
        x"2D0E",
        x"2D1F",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"239E",
        x"0F99",
        x"0B66",
        x"2F76",
        x"2F86",
        x"2F97",
        x"940E",
        x"22C6",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"22B2",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"1BCA",
        x"0BDB",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"9409",
        x"882A",
        x"8839",
        x"8848",
        x"845F",
        x"846E",
        x"847D",
        x"848C",
        x"849B",
        x"84AA",
        x"84B9",
        x"84C8",
        x"80DF",
        x"80EE",
        x"80FD",
        x"810C",
        x"811B",
        x"81AA",
        x"81B9",
        x"0FCE",
        x"1DD1",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2FCA",
        x"2FDB",
        x"9508",
        x"93DF",
        x"93CF",
        x"929F",
        x"E4A0",
        x"2E9A",
        x"2400",
        x"2DA0",
        x"2DB1",
        x"2DC0",
        x"2DD1",
        x"2DE0",
        x"2DF1",
        x"9516",
        x"9507",
        x"94F7",
        x"94E7",
        x"94D7",
        x"94C7",
        x"94B7",
        x"94A7",
        x"F448",
        x"6810",
        x"0FA2",
        x"1FB3",
        x"1FC4",
        x"1FD5",
        x"1FE6",
        x"1FF7",
        x"1E08",
        x"1E19",
        x"0F22",
        x"1F33",
        x"1F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"949A",
        x"F721",
        x"2F2A",
        x"2F3B",
        x"2F4C",
        x"2F5D",
        x"2F6E",
        x"2F7F",
        x"2D80",
        x"2D91",
        x"2411",
        x"909F",
        x"91CF",
        x"91DF",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"95C8",
        x"9631",
        x"920D",
        x"2000",
        x"F7D9",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"5041",
        x"4050",
        x"F050",
        x"95C8",
        x"9631",
        x"920D",
        x"2000",
        x"F7C1",
        x"C001",
        x"921D",
        x"5041",
        x"4050",
        x"F7E0",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"C004",
        x"918D",
        x"9001",
        x"1980",
        x"F421",
        x"5041",
        x"4050",
        x"F7C8",
        x"1B88",
        x"0B99",
        x"9508",
        x"2FA8",
        x"2FB9",
        x"C001",
        x"936D",
        x"5041",
        x"4050",
        x"F7E0",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"9001",
        x"920D",
        x"2000",
        x"F7E1",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"5041",
        x"4050",
        x"F048",
        x"9001",
        x"920D",
        x"2000",
        x"F7C9",
        x"C001",
        x"921D",
        x"5041",
        x"4050",
        x"F7E0",
        x"9508",
        x"99E1",
        x"CFFE",
        x"BB9F",
        x"BB8E",
        x"9AE0",
        x"2799",
        x"B38D",
        x"9508",
        x"2F26",
        x"99E1",
        x"CFFE",
        x"BB9F",
        x"BB8E",
        x"BB2D",
        x"B60F",
        x"94F8",
        x"9AE2",
        x"9AE1",
        x"BE0F",
        x"9601",
        x"9508",
        x"94F8",
        x"CFFF",
        x"FF55",
        x"FFFF",
        x"18FF",
        x"E921",
        x"DE20",
        x"7B20",
        x"1720",
        x"C820",
        x"7A1F",
        x"511F",
        x"C221",
        x"B51E",
        x"A01E",
        x"6C1E",
        x"211E",
        x"AF1E",
        x"A31D",
        x"971D",
        x"781D",
        x"641D",
        x"571D",
        x"4A1D",
        x"3D1D",
        x"CA1D",
        x"AF1C",
        x"201C",
        x"2A22",
        x"2C2B",
        x"3D5B",
        x"7C5D",
        x"007F",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000"
    );

begin

    process (cp2)
    begin
        if rising_edge(cp2) then
            if ce = '1' then
                if (we = '1') then
                    RAM(conv_integer(address)) <= din;
                end if;
                dout <= RAM(conv_integer(address));
            end if;
        end if;
    end process;

end RTL;

