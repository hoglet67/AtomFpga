library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mc6847_ntsc is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of mc6847_ntsc is

  signal rom_addr : std_logic_vector(9 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(9 downto 0) <= ADDR(9 downto 0);
  end process;

  p_rom : process
  begin
    wait until rising_edge(CLK);
    DATA <= (others => '0');
  
 if  rom_addr(9 downto 8) = "00" then
	 case rom_addr(7 downto 0) is
      when x"00" => DATA <= x"00";
      when x"01" => DATA <= x"00";
      when x"02" => DATA <= x"00";
      when x"03" => DATA <= x"1C";
      when x"04" => DATA <= x"22";
      when x"05" => DATA <= x"02";
      when x"06" => DATA <= x"1A";
      when x"07" => DATA <= x"2A";
      when x"08" => DATA <= x"2A";
      when x"09" => DATA <= x"1C";
      when x"0A" => DATA <= x"00";
      when x"0B" => DATA <= x"00";
		when x"0C" => DATA <= x"00";
      when x"0D" => DATA <= x"00";
      when x"0E" => DATA <= x"00";
      when x"0F" => DATA <= x"00";
		when x"10" => DATA <= x"00";
      when x"11" => DATA <= x"00";
      when x"12" => DATA <= x"00";
      when x"13" => DATA <= x"08";
      when x"14" => DATA <= x"14";
      when x"15" => DATA <= x"22";
      when x"16" => DATA <= x"22";
      when x"17" => DATA <= x"3E";
      when x"18" => DATA <= x"22";
      when x"19" => DATA <= x"22";
      when x"1A" => DATA <= x"00";
      when x"1B" => DATA <= x"00";
      when x"1C" => DATA <= x"00";
      when x"1D" => DATA <= x"00";
      when x"1E" => DATA <= x"00";
      when x"1F" => DATA <= x"00";
      when x"20" => DATA <= x"00";
      when x"21" => DATA <= x"00";
      when x"22" => DATA <= x"00";
      when x"23" => DATA <= x"3C";
      when x"24" => DATA <= x"12";
      when x"25" => DATA <= x"12";
      when x"26" => DATA <= x"1C";
      when x"27" => DATA <= x"12";
      when x"28" => DATA <= x"12";
      when x"29" => DATA <= x"3C";
      when x"2A" => DATA <= x"00";
      when x"2B" => DATA <= x"00";
      when x"2C" => DATA <= x"00";
      when x"2D" => DATA <= x"00";
      when x"2E" => DATA <= x"00";
      when x"2F" => DATA <= x"00";
      when x"30" => DATA <= x"00";
      when x"31" => DATA <= x"00";
      when x"32" => DATA <= x"00";
      when x"33" => DATA <= x"1C";
      when x"34" => DATA <= x"22";
      when x"35" => DATA <= x"20";
      when x"36" => DATA <= x"20";
      when x"37" => DATA <= x"20";
      when x"38" => DATA <= x"22";
      when x"39" => DATA <= x"1C";
      when x"3A" => DATA <= x"00";
      when x"3B" => DATA <= x"00";
      when x"3C" => DATA <= x"00";
      when x"3D" => DATA <= x"00";
      when x"3E" => DATA <= x"00";
      when x"3F" => DATA <= x"00";
      when x"40" => DATA <= x"00";
      when x"41" => DATA <= x"00";
      when x"42" => DATA <= x"00";
      when x"43" => DATA <= x"3C";
      when x"44" => DATA <= x"12";
      when x"45" => DATA <= x"12";
      when x"46" => DATA <= x"12";
      when x"47" => DATA <= x"12";
      when x"48" => DATA <= x"12";
      when x"49" => DATA <= x"3C";
      when x"4A" => DATA <= x"00";
      when x"4B" => DATA <= x"00";
      when x"4C" => DATA <= x"00";
      when x"4D" => DATA <= x"00";
      when x"4E" => DATA <= x"00";
      when x"4F" => DATA <= x"00";
      when x"50" => DATA <= x"00";
      when x"51" => DATA <= x"00";
      when x"52" => DATA <= x"00";
      when x"53" => DATA <= x"3E";
      when x"54" => DATA <= x"20";
      when x"55" => DATA <= x"20";
      when x"56" => DATA <= x"38";
      when x"57" => DATA <= x"20";
      when x"58" => DATA <= x"20";
      when x"59" => DATA <= x"3E";
      when x"5A" => DATA <= x"00";
      when x"5B" => DATA <= x"00";
      when x"5C" => DATA <= x"00";
      when x"5D" => DATA <= x"00";
      when x"5E" => DATA <= x"00";
      when x"5F" => DATA <= x"00";
      when x"60" => DATA <= x"00";
      when x"61" => DATA <= x"00";
      when x"62" => DATA <= x"00";
      when x"63" => DATA <= x"3E";
      when x"64" => DATA <= x"20";
      when x"65" => DATA <= x"20";
      when x"66" => DATA <= x"38";
      when x"67" => DATA <= x"20";
      when x"68" => DATA <= x"20";
      when x"69" => DATA <= x"20";
      when x"6A" => DATA <= x"00";
      when x"6B" => DATA <= x"00";
      when x"6C" => DATA <= x"00";
      when x"6D" => DATA <= x"00";
      when x"6E" => DATA <= x"00";
      when x"6F" => DATA <= x"00";
      when x"70" => DATA <= x"00";
      when x"71" => DATA <= x"00";
      when x"72" => DATA <= x"00";
      when x"73" => DATA <= x"1E";
      when x"74" => DATA <= x"20";
      when x"75" => DATA <= x"20";
      when x"76" => DATA <= x"26";
      when x"77" => DATA <= x"22";
      when x"78" => DATA <= x"22";
      when x"79" => DATA <= x"1E";
      when x"7A" => DATA <= x"00";
      when x"7B" => DATA <= x"00";
      when x"7C" => DATA <= x"00";
      when x"7D" => DATA <= x"00";
      when x"7E" => DATA <= x"00";
      when x"7F" => DATA <= x"00";
      when x"80" => DATA <= x"00";
      when x"81" => DATA <= x"00";
      when x"82" => DATA <= x"00";
      when x"83" => DATA <= x"22";
      when x"84" => DATA <= x"22";
      when x"85" => DATA <= x"22";
      when x"86" => DATA <= x"3E";
      when x"87" => DATA <= x"22";
      when x"88" => DATA <= x"22";
      when x"89" => DATA <= x"22";
      when x"8A" => DATA <= x"00";
      when x"8B" => DATA <= x"00";
      when x"8C" => DATA <= x"00";
      when x"8D" => DATA <= x"00";
      when x"8E" => DATA <= x"00";
      when x"8F" => DATA <= x"00";
      when x"90" => DATA <= x"00";
      when x"91" => DATA <= x"00";
      when x"92" => DATA <= x"00";
      when x"93" => DATA <= x"1C";
      when x"94" => DATA <= x"08";
      when x"95" => DATA <= x"08";
      when x"96" => DATA <= x"08";
      when x"97" => DATA <= x"08";
      when x"98" => DATA <= x"08";
      when x"99" => DATA <= x"1C";
      when x"9A" => DATA <= x"00";
      when x"9B" => DATA <= x"00";
      when x"9C" => DATA <= x"00";
      when x"9D" => DATA <= x"00";
      when x"9E" => DATA <= x"00";
      when x"9F" => DATA <= x"00";
      when x"A0" => DATA <= x"00";
      when x"A1" => DATA <= x"00";
      when x"A2" => DATA <= x"00";
      when x"A3" => DATA <= x"02";
      when x"A4" => DATA <= x"02";
      when x"A5" => DATA <= x"02";
      when x"A6" => DATA <= x"02";
      when x"A7" => DATA <= x"22";
      when x"A8" => DATA <= x"22";
      when x"A9" => DATA <= x"1C";
      when x"AA" => DATA <= x"00";
      when x"AB" => DATA <= x"00";
      when x"AC" => DATA <= x"00";
      when x"AD" => DATA <= x"00";
      when x"AE" => DATA <= x"00";
      when x"AF" => DATA <= x"00";
      when x"B0" => DATA <= x"00";
      when x"B1" => DATA <= x"00";
      when x"B2" => DATA <= x"00";
      when x"B3" => DATA <= x"22";
      when x"B4" => DATA <= x"24";
      when x"B5" => DATA <= x"28";
      when x"B6" => DATA <= x"30";
      when x"B7" => DATA <= x"28";
      when x"B8" => DATA <= x"24";
      when x"B9" => DATA <= x"22";
      when x"BA" => DATA <= x"00";
      when x"BB" => DATA <= x"00";
      when x"BC" => DATA <= x"00";
      when x"BD" => DATA <= x"00";
      when x"BE" => DATA <= x"00";
      when x"BF" => DATA <= x"00";
      when x"C0" => DATA <= x"00";
      when x"C1" => DATA <= x"00";
      when x"C2" => DATA <= x"00";
      when x"C3" => DATA <= x"20";
      when x"C4" => DATA <= x"20";
      when x"C5" => DATA <= x"20";
      when x"C6" => DATA <= x"20";
      when x"C7" => DATA <= x"20";
      when x"C8" => DATA <= x"20";
      when x"C9" => DATA <= x"3E";
      when x"CA" => DATA <= x"00";
      when x"CB" => DATA <= x"00";
      when x"CC" => DATA <= x"00";
      when x"CD" => DATA <= x"00";
      when x"CE" => DATA <= x"00";
      when x"CF" => DATA <= x"00";
      when x"D0" => DATA <= x"00";
      when x"D1" => DATA <= x"00";
      when x"D2" => DATA <= x"00";
      when x"D3" => DATA <= x"22";
      when x"D4" => DATA <= x"36";
      when x"D5" => DATA <= x"2A";
      when x"D6" => DATA <= x"2A";
      when x"D7" => DATA <= x"22";
      when x"D8" => DATA <= x"22";
      when x"D9" => DATA <= x"22";
      when x"DA" => DATA <= x"00";
      when x"DB" => DATA <= x"00";
      when x"DC" => DATA <= x"00";
      when x"DD" => DATA <= x"00";
      when x"DE" => DATA <= x"00";
      when x"DF" => DATA <= x"00";
      when x"E0" => DATA <= x"00";
      when x"E1" => DATA <= x"00";
      when x"E2" => DATA <= x"00";
      when x"E3" => DATA <= x"22";
      when x"E4" => DATA <= x"32";
      when x"E5" => DATA <= x"2A";
      when x"E6" => DATA <= x"26";
      when x"E7" => DATA <= x"22";
      when x"E8" => DATA <= x"22";
      when x"E9" => DATA <= x"22";
      when x"EA" => DATA <= x"00";
      when x"EB" => DATA <= x"00";
      when x"EC" => DATA <= x"00";
      when x"ED" => DATA <= x"00";
      when x"EE" => DATA <= x"00";
      when x"EF" => DATA <= x"00";
      when x"F0" => DATA <= x"00";
      when x"F1" => DATA <= x"00";
      when x"F2" => DATA <= x"00";
      when x"F3" => DATA <= x"3E";
      when x"F4" => DATA <= x"22";
      when x"F5" => DATA <= x"22";
      when x"F6" => DATA <= x"22";
      when x"F7" => DATA <= x"22";
      when x"F8" => DATA <= x"22";
      when x"F9" => DATA <= x"3E";
      when x"FA" => DATA <= x"00";
      when x"FB" => DATA <= x"00";
      when x"FC" => DATA <= x"00";
      when x"FD" => DATA <= x"00";
      when x"FE" => DATA <= x"00";
      when x"FF" => DATA <= x"00";
		when others => DATA <= (others => '0');
    end case;
end if;	


if  rom_addr(9 downto 8) = "01" then	
   case rom_addr(7 downto 0) is
      when x"00" => DATA <= x"00";
      when x"01" => DATA <= x"00";
      when x"02" => DATA <= x"00";
      when x"03" => DATA <= x"3C";
      when x"04" => DATA <= x"22";
      when x"05" => DATA <= x"22";
      when x"06" => DATA <= x"3C";
      when x"07" => DATA <= x"20";
      when x"08" => DATA <= x"20";
      when x"09" => DATA <= x"20";
      when x"0A" => DATA <= x"00";
      when x"0B" => DATA <= x"00";
      when x"0C" => DATA <= x"00";
      when x"0D" => DATA <= x"00";
      when x"0E" => DATA <= x"00";
      when x"0F" => DATA <= x"00";
      when x"10" => DATA <= x"00";
      when x"11" => DATA <= x"00";
      when x"12" => DATA <= x"00";
      when x"13" => DATA <= x"1C";
      when x"14" => DATA <= x"22";
      when x"15" => DATA <= x"22";
      when x"16" => DATA <= x"22";
      when x"17" => DATA <= x"2A";
      when x"18" => DATA <= x"24";
      when x"19" => DATA <= x"1A";
      when x"1A" => DATA <= x"00";
      when x"1B" => DATA <= x"00";
      when x"1C" => DATA <= x"00";
      when x"1D" => DATA <= x"00";
      when x"1E" => DATA <= x"00";
      when x"1F" => DATA <= x"00";
      when x"20" => DATA <= x"00";
      when x"21" => DATA <= x"00";
      when x"22" => DATA <= x"00";
      when x"23" => DATA <= x"3C";
      when x"24" => DATA <= x"22";
      when x"25" => DATA <= x"22";
      when x"26" => DATA <= x"3C";
      when x"27" => DATA <= x"28";
      when x"28" => DATA <= x"24";
      when x"29" => DATA <= x"22";
      when x"2A" => DATA <= x"00";
      when x"2B" => DATA <= x"00";
      when x"2C" => DATA <= x"00";
      when x"2D" => DATA <= x"00";
      when x"2E" => DATA <= x"00";
      when x"2F" => DATA <= x"00";
      when x"30" => DATA <= x"00";
      when x"31" => DATA <= x"00";
      when x"32" => DATA <= x"00";
      when x"33" => DATA <= x"1C";
      when x"34" => DATA <= x"22";
      when x"35" => DATA <= x"10";
      when x"36" => DATA <= x"08";
      when x"37" => DATA <= x"04";
      when x"38" => DATA <= x"22";
      when x"39" => DATA <= x"1C";
      when x"3A" => DATA <= x"00";
      when x"3B" => DATA <= x"00";
      when x"3C" => DATA <= x"00";
      when x"3D" => DATA <= x"00";
      when x"3E" => DATA <= x"00";
      when x"3F" => DATA <= x"00";
      when x"40" => DATA <= x"00";
      when x"41" => DATA <= x"00";
      when x"42" => DATA <= x"00";
      when x"43" => DATA <= x"3E";
      when x"44" => DATA <= x"08";
      when x"45" => DATA <= x"08";
      when x"46" => DATA <= x"08";
      when x"47" => DATA <= x"08";
      when x"48" => DATA <= x"08";
      when x"49" => DATA <= x"08";
      when x"4A" => DATA <= x"00";
      when x"4B" => DATA <= x"00";
      when x"4C" => DATA <= x"00";
      when x"4D" => DATA <= x"00";
      when x"4E" => DATA <= x"00";
      when x"4F" => DATA <= x"00";
      when x"50" => DATA <= x"00";
      when x"51" => DATA <= x"00";
      when x"52" => DATA <= x"00";
      when x"53" => DATA <= x"22";
      when x"54" => DATA <= x"22";
      when x"55" => DATA <= x"22";
      when x"56" => DATA <= x"22";
      when x"57" => DATA <= x"22";
      when x"58" => DATA <= x"22";
      when x"59" => DATA <= x"1C";
      when x"5A" => DATA <= x"00";
      when x"5B" => DATA <= x"00";
      when x"5C" => DATA <= x"00";
      when x"5D" => DATA <= x"00";
      when x"5E" => DATA <= x"00";
      when x"5F" => DATA <= x"00";
      when x"60" => DATA <= x"00";
      when x"61" => DATA <= x"00";
      when x"62" => DATA <= x"00";
      when x"63" => DATA <= x"22";
      when x"64" => DATA <= x"22";
      when x"65" => DATA <= x"22";
      when x"66" => DATA <= x"14";
      when x"67" => DATA <= x"14";
      when x"68" => DATA <= x"08";
      when x"69" => DATA <= x"08";
      when x"6A" => DATA <= x"00";
      when x"6B" => DATA <= x"00";
      when x"6C" => DATA <= x"00";
      when x"6D" => DATA <= x"00";
      when x"6E" => DATA <= x"00";
      when x"6F" => DATA <= x"00";
      when x"70" => DATA <= x"00";
      when x"71" => DATA <= x"00";
      when x"72" => DATA <= x"00";
      when x"73" => DATA <= x"22";
      when x"74" => DATA <= x"22";
      when x"75" => DATA <= x"22";
      when x"76" => DATA <= x"2A";
      when x"77" => DATA <= x"2A";
      when x"78" => DATA <= x"36";
      when x"79" => DATA <= x"22";
      when x"7A" => DATA <= x"00";
      when x"7B" => DATA <= x"00";
      when x"7C" => DATA <= x"00";
      when x"7D" => DATA <= x"00";
      when x"7E" => DATA <= x"00";
      when x"7F" => DATA <= x"00";
      when x"80" => DATA <= x"00";
      when x"81" => DATA <= x"00";
      when x"82" => DATA <= x"00";
      when x"83" => DATA <= x"22";
      when x"84" => DATA <= x"22";
      when x"85" => DATA <= x"14";
      when x"86" => DATA <= x"08";
      when x"87" => DATA <= x"14";
      when x"88" => DATA <= x"22";
      when x"89" => DATA <= x"22";
      when x"8A" => DATA <= x"00";
      when x"8B" => DATA <= x"00";
      when x"8C" => DATA <= x"00";
      when x"8D" => DATA <= x"00";
      when x"8E" => DATA <= x"00";
      when x"8F" => DATA <= x"00";
      when x"90" => DATA <= x"00";
      when x"91" => DATA <= x"00";
      when x"92" => DATA <= x"00";
      when x"93" => DATA <= x"22";
      when x"94" => DATA <= x"22";
      when x"95" => DATA <= x"14";
      when x"96" => DATA <= x"08";
      when x"97" => DATA <= x"08";
      when x"98" => DATA <= x"08";
      when x"99" => DATA <= x"08";
      when x"9A" => DATA <= x"00";
      when x"9B" => DATA <= x"00";
      when x"9C" => DATA <= x"00";
      when x"9D" => DATA <= x"00";
      when x"9E" => DATA <= x"00";
      when x"9F" => DATA <= x"00";
      when x"A0" => DATA <= x"00";
      when x"A1" => DATA <= x"00";
      when x"A2" => DATA <= x"00";
      when x"A3" => DATA <= x"3E";
      when x"A4" => DATA <= x"02";
      when x"A5" => DATA <= x"04";
      when x"A6" => DATA <= x"08";
      when x"A7" => DATA <= x"10";
      when x"A8" => DATA <= x"20";
      when x"A9" => DATA <= x"3E";
      when x"AA" => DATA <= x"00";
      when x"AB" => DATA <= x"00";
      when x"AC" => DATA <= x"00";
      when x"AD" => DATA <= x"00";
      when x"AE" => DATA <= x"00";
      when x"AF" => DATA <= x"00";
      when x"B0" => DATA <= x"00";
      when x"B1" => DATA <= x"00";
      when x"B2" => DATA <= x"00";
      when x"B3" => DATA <= x"38";
      when x"B4" => DATA <= x"20";
      when x"B5" => DATA <= x"20";
      when x"B6" => DATA <= x"20";
      when x"B7" => DATA <= x"20";
      when x"B8" => DATA <= x"20";
      when x"B9" => DATA <= x"38";
      when x"BA" => DATA <= x"00";
      when x"BB" => DATA <= x"00";
      when x"BC" => DATA <= x"00";
      when x"BD" => DATA <= x"00";
      when x"BE" => DATA <= x"00";
      when x"BF" => DATA <= x"00";
      when x"C0" => DATA <= x"00";
      when x"C1" => DATA <= x"00";
      when x"C2" => DATA <= x"00";
      when x"C3" => DATA <= x"20";
      when x"C4" => DATA <= x"20";
      when x"C5" => DATA <= x"10";
      when x"C6" => DATA <= x"08";
      when x"C7" => DATA <= x"04";
      when x"C8" => DATA <= x"02";
      when x"C9" => DATA <= x"02";
      when x"CA" => DATA <= x"00";
      when x"CB" => DATA <= x"00";
      when x"CC" => DATA <= x"00";
      when x"CD" => DATA <= x"00";
      when x"CE" => DATA <= x"00";
      when x"CF" => DATA <= x"00";
      when x"D0" => DATA <= x"00";
      when x"D1" => DATA <= x"00";
      when x"D2" => DATA <= x"00";
      when x"D3" => DATA <= x"0E";
      when x"D4" => DATA <= x"02";
      when x"D5" => DATA <= x"02";
      when x"D6" => DATA <= x"02";
      when x"D7" => DATA <= x"02";
      when x"D8" => DATA <= x"02";
      when x"D9" => DATA <= x"0E";
      when x"DA" => DATA <= x"00";
      when x"DB" => DATA <= x"00";
      when x"DC" => DATA <= x"00";
      when x"DD" => DATA <= x"00";
      when x"DE" => DATA <= x"00";
      when x"DF" => DATA <= x"00";
      when x"E0" => DATA <= x"00";
      when x"E1" => DATA <= x"00";
      when x"E2" => DATA <= x"00";
      when x"E3" => DATA <= x"08";
      when x"E4" => DATA <= x"1C";
      when x"E5" => DATA <= x"2A";
      when x"E6" => DATA <= x"08";
      when x"E7" => DATA <= x"08";
      when x"E8" => DATA <= x"08";
      when x"E9" => DATA <= x"08";
      when x"EA" => DATA <= x"00";
      when x"EB" => DATA <= x"00";
      when x"EC" => DATA <= x"00";
      when x"ED" => DATA <= x"00";
      when x"EE" => DATA <= x"00";
      when x"EF" => DATA <= x"00";
      when x"F0" => DATA <= x"00";
      when x"F1" => DATA <= x"00";
      when x"F2" => DATA <= x"00";
      when x"F3" => DATA <= x"00";
      when x"F4" => DATA <= x"08";
      when x"F5" => DATA <= x"10";
      when x"F6" => DATA <= x"3E";
      when x"F7" => DATA <= x"10";
      when x"F8" => DATA <= x"08";
      when x"F9" => DATA <= x"00";
      when x"FA" => DATA <= x"00";
      when x"FB" => DATA <= x"00";
      when x"FC" => DATA <= x"00";
      when x"FD" => DATA <= x"00";
      when x"FE" => DATA <= x"00";
      when x"FF" => DATA <= x"00";
      when others => DATA <= (others => '0');
	   end case;
end if;	


if  rom_addr(9 downto 8) = "10" then	
   case rom_addr(7 downto 0) is
	  when x"00" => DATA <= x"00";
      when x"01" => DATA <= x"00";
      when x"02" => DATA <= x"00";
      when x"03" => DATA <= x"00";
      when x"04" => DATA <= x"00";
      when x"05" => DATA <= x"00";
      when x"06" => DATA <= x"00";
      when x"07" => DATA <= x"00";
      when x"08" => DATA <= x"00";
      when x"09" => DATA <= x"00";
      when x"0A" => DATA <= x"00";
      when x"0B" => DATA <= x"00";
      when x"0C" => DATA <= x"00";
      when x"0D" => DATA <= x"00";
      when x"0E" => DATA <= x"00";
      when x"0F" => DATA <= x"00";
      when x"10" => DATA <= x"00";
      when x"11" => DATA <= x"00";
      when x"12" => DATA <= x"00";
      when x"13" => DATA <= x"08";
      when x"14" => DATA <= x"08";
      when x"15" => DATA <= x"08";
      when x"16" => DATA <= x"08";
      when x"17" => DATA <= x"08";
      when x"18" => DATA <= x"00";
      when x"19" => DATA <= x"08";
      when x"1A" => DATA <= x"00";
      when x"1B" => DATA <= x"00";
      when x"1C" => DATA <= x"00";
      when x"1D" => DATA <= x"00";
      when x"1E" => DATA <= x"00";
      when x"1F" => DATA <= x"00";
      when x"20" => DATA <= x"00";
      when x"21" => DATA <= x"00";
      when x"22" => DATA <= x"00";
      when x"23" => DATA <= x"14";
      when x"24" => DATA <= x"14";
      when x"25" => DATA <= x"14";
      when x"26" => DATA <= x"00";
      when x"27" => DATA <= x"00";
      when x"28" => DATA <= x"00";
      when x"29" => DATA <= x"00";
      when x"2A" => DATA <= x"00";
      when x"2B" => DATA <= x"00";
      when x"2C" => DATA <= x"00";
      when x"2D" => DATA <= x"00";
      when x"2E" => DATA <= x"00";
      when x"2F" => DATA <= x"00";
      when x"30" => DATA <= x"00";
      when x"31" => DATA <= x"00";
      when x"32" => DATA <= x"00";
      when x"33" => DATA <= x"14";
      when x"34" => DATA <= x"14";
      when x"35" => DATA <= x"36";
      when x"36" => DATA <= x"00";
      when x"37" => DATA <= x"36";
      when x"38" => DATA <= x"14";
      when x"39" => DATA <= x"14";
      when x"3A" => DATA <= x"00";
      when x"3B" => DATA <= x"00";
      when x"3C" => DATA <= x"00";
      when x"3D" => DATA <= x"00";
      when x"3E" => DATA <= x"00";
      when x"3F" => DATA <= x"00";
      when x"40" => DATA <= x"00";
      when x"41" => DATA <= x"00";
      when x"42" => DATA <= x"00";
      when x"43" => DATA <= x"08";
      when x"44" => DATA <= x"1E";
      when x"45" => DATA <= x"20";
      when x"46" => DATA <= x"1C";
      when x"47" => DATA <= x"02";
      when x"48" => DATA <= x"3C";
      when x"49" => DATA <= x"08";
      when x"4A" => DATA <= x"00";
      when x"4B" => DATA <= x"00";
      when x"4C" => DATA <= x"00";
      when x"4D" => DATA <= x"00";
      when x"4E" => DATA <= x"00";
      when x"4F" => DATA <= x"00";
      when x"50" => DATA <= x"00";
      when x"51" => DATA <= x"00";
      when x"52" => DATA <= x"00";
      when x"53" => DATA <= x"32";
      when x"54" => DATA <= x"32";
      when x"55" => DATA <= x"04";
      when x"56" => DATA <= x"08";
      when x"57" => DATA <= x"10";
      when x"58" => DATA <= x"26";
      when x"59" => DATA <= x"26";
      when x"5A" => DATA <= x"00";
      when x"5B" => DATA <= x"00";
      when x"5C" => DATA <= x"00";
      when x"5D" => DATA <= x"00";
      when x"5E" => DATA <= x"00";
      when x"5F" => DATA <= x"00";
      when x"60" => DATA <= x"00";
      when x"61" => DATA <= x"00";
      when x"62" => DATA <= x"00";
      when x"63" => DATA <= x"10";
      when x"64" => DATA <= x"28";
      when x"65" => DATA <= x"28";
      when x"66" => DATA <= x"10";
      when x"67" => DATA <= x"2A";
      when x"68" => DATA <= x"24";
      when x"69" => DATA <= x"1A";
      when x"6A" => DATA <= x"00";
      when x"6B" => DATA <= x"00";
      when x"6C" => DATA <= x"00";
      when x"6D" => DATA <= x"00";
      when x"6E" => DATA <= x"00";
      when x"6F" => DATA <= x"00";
      when x"70" => DATA <= x"00";
      when x"71" => DATA <= x"00";
      when x"72" => DATA <= x"00";
      when x"73" => DATA <= x"18";
      when x"74" => DATA <= x"18";
      when x"75" => DATA <= x"18";
      when x"76" => DATA <= x"00";
      when x"77" => DATA <= x"00";
      when x"78" => DATA <= x"00";
      when x"79" => DATA <= x"00";
      when x"7A" => DATA <= x"00";
      when x"7B" => DATA <= x"00";
      when x"7C" => DATA <= x"00";
      when x"7D" => DATA <= x"00";
      when x"7E" => DATA <= x"00";
      when x"7F" => DATA <= x"00";
      when x"80" => DATA <= x"00";
      when x"81" => DATA <= x"00";
      when x"82" => DATA <= x"00";
      when x"83" => DATA <= x"08";
      when x"84" => DATA <= x"10";
      when x"85" => DATA <= x"20";
      when x"86" => DATA <= x"20";
      when x"87" => DATA <= x"20";
      when x"88" => DATA <= x"10";
      when x"89" => DATA <= x"08";
      when x"8A" => DATA <= x"00";
      when x"8B" => DATA <= x"00";
      when x"8C" => DATA <= x"00";
      when x"8D" => DATA <= x"00";
      when x"8E" => DATA <= x"00";
      when x"8F" => DATA <= x"00";
      when x"90" => DATA <= x"00";
      when x"91" => DATA <= x"00";
      when x"92" => DATA <= x"00";
      when x"93" => DATA <= x"08";
      when x"94" => DATA <= x"04";
      when x"95" => DATA <= x"02";
      when x"96" => DATA <= x"02";
      when x"97" => DATA <= x"02";
      when x"98" => DATA <= x"04";
      when x"99" => DATA <= x"08";
      when x"9A" => DATA <= x"00";
      when x"9B" => DATA <= x"00";
      when x"9C" => DATA <= x"00";
      when x"9D" => DATA <= x"00";
      when x"9E" => DATA <= x"00";
      when x"9F" => DATA <= x"00";
      when x"A0" => DATA <= x"00";
      when x"A1" => DATA <= x"00";
      when x"A2" => DATA <= x"00";
      when x"A3" => DATA <= x"00";
      when x"A4" => DATA <= x"08";
      when x"A5" => DATA <= x"1C";
      when x"A6" => DATA <= x"3E";
      when x"A7" => DATA <= x"1C";
      when x"A8" => DATA <= x"08";
      when x"A9" => DATA <= x"00";
      when x"AA" => DATA <= x"00";
      when x"AB" => DATA <= x"00";
      when x"AC" => DATA <= x"00";
      when x"AD" => DATA <= x"00";
      when x"AE" => DATA <= x"00";
      when x"AF" => DATA <= x"00";
      when x"B0" => DATA <= x"00";
      when x"B1" => DATA <= x"00";
      when x"B2" => DATA <= x"00";
      when x"B3" => DATA <= x"00";
      when x"B4" => DATA <= x"08";
      when x"B5" => DATA <= x"08";
      when x"B6" => DATA <= x"3E";
      when x"B7" => DATA <= x"08";
      when x"B8" => DATA <= x"08";
      when x"B9" => DATA <= x"00";
      when x"BA" => DATA <= x"00";
      when x"BB" => DATA <= x"00";
      when x"BC" => DATA <= x"00";
      when x"BD" => DATA <= x"00";
      when x"BE" => DATA <= x"00";
      when x"BF" => DATA <= x"00";
      when x"C0" => DATA <= x"00";
      when x"C1" => DATA <= x"00";
      when x"C2" => DATA <= x"00";
      when x"C3" => DATA <= x"00";
      when x"C4" => DATA <= x"00";
      when x"C5" => DATA <= x"00";
      when x"C6" => DATA <= x"30";
      when x"C7" => DATA <= x"30";
      when x"C8" => DATA <= x"10";
      when x"C9" => DATA <= x"20";
      when x"CA" => DATA <= x"00";
      when x"CB" => DATA <= x"00";
      when x"CC" => DATA <= x"00";
      when x"CD" => DATA <= x"00";
      when x"CE" => DATA <= x"00";
      when x"CF" => DATA <= x"00";
      when x"D0" => DATA <= x"00";
      when x"D1" => DATA <= x"00";
      when x"D2" => DATA <= x"00";
      when x"D3" => DATA <= x"00";
      when x"D4" => DATA <= x"00";
      when x"D5" => DATA <= x"00";
      when x"D6" => DATA <= x"3E";
      when x"D7" => DATA <= x"00";
      when x"D8" => DATA <= x"00";
      when x"D9" => DATA <= x"00";
      when x"DA" => DATA <= x"00";
      when x"DB" => DATA <= x"00";
      when x"DC" => DATA <= x"00";
      when x"DD" => DATA <= x"00";
      when x"DE" => DATA <= x"00";
      when x"DF" => DATA <= x"00";
      when x"E0" => DATA <= x"00";
      when x"E1" => DATA <= x"00";
      when x"E2" => DATA <= x"00";
      when x"E3" => DATA <= x"00";
      when x"E4" => DATA <= x"00";
      when x"E5" => DATA <= x"00";
      when x"E6" => DATA <= x"00";
      when x"E7" => DATA <= x"00";
      when x"E8" => DATA <= x"30";
      when x"E9" => DATA <= x"30";
      when x"EA" => DATA <= x"00";
      when x"EB" => DATA <= x"00";
      when x"EC" => DATA <= x"00";
      when x"ED" => DATA <= x"00";
      when x"EE" => DATA <= x"00";
      when x"EF" => DATA <= x"00";
      when x"F0" => DATA <= x"00";
      when x"F1" => DATA <= x"00";
      when x"F2" => DATA <= x"00";
      when x"F3" => DATA <= x"02";
      when x"F4" => DATA <= x"02";
      when x"F5" => DATA <= x"04";
      when x"F6" => DATA <= x"08";
      when x"F7" => DATA <= x"10";
      when x"F8" => DATA <= x"20";
      when x"F9" => DATA <= x"20";
      when x"FA" => DATA <= x"00";
      when x"FB" => DATA <= x"00";
      when x"FC" => DATA <= x"00";
      when x"FD" => DATA <= x"00";
      when x"FE" => DATA <= x"00";
      when x"FF" => DATA <= x"00";
		when others => DATA <= (others => '0');
	   end case;
end if;	


if  rom_addr(9 downto 8) = "11" then	
   case rom_addr(7 downto 0) is		
     when x"00" => DATA <= x"00";
      when x"01" => DATA <= x"00";
      when x"02" => DATA <= x"00";
      when x"03" => DATA <= x"18";
      when x"04" => DATA <= x"24";
      when x"05" => DATA <= x"24";
      when x"06" => DATA <= x"24";
      when x"07" => DATA <= x"24";
      when x"08" => DATA <= x"24";
      when x"09" => DATA <= x"18";
      when x"0A" => DATA <= x"00";
      when x"0B" => DATA <= x"00";
      when x"0C" => DATA <= x"00";
      when x"0D" => DATA <= x"00";
      when x"0E" => DATA <= x"00";
      when x"0F" => DATA <= x"00";
      when x"10" => DATA <= x"00";
      when x"11" => DATA <= x"00";
      when x"12" => DATA <= x"00";
      when x"13" => DATA <= x"08";
      when x"14" => DATA <= x"18";
      when x"15" => DATA <= x"08";
      when x"16" => DATA <= x"08";
      when x"17" => DATA <= x"08";
      when x"18" => DATA <= x"08";
      when x"19" => DATA <= x"1C";
      when x"1A" => DATA <= x"00";
      when x"1B" => DATA <= x"00";
      when x"1C" => DATA <= x"00";
      when x"1D" => DATA <= x"00";
      when x"1E" => DATA <= x"00";
      when x"1F" => DATA <= x"00";
      when x"20" => DATA <= x"00";
      when x"21" => DATA <= x"00";
      when x"22" => DATA <= x"00";
      when x"23" => DATA <= x"1C";
      when x"24" => DATA <= x"22";
      when x"25" => DATA <= x"02";
      when x"26" => DATA <= x"1C";
      when x"27" => DATA <= x"20";
      when x"28" => DATA <= x"20";
      when x"29" => DATA <= x"3E";
      when x"2A" => DATA <= x"00";
      when x"2B" => DATA <= x"00";
      when x"2C" => DATA <= x"00";
      when x"2D" => DATA <= x"00";
      when x"2E" => DATA <= x"00";
      when x"2F" => DATA <= x"00";
      when x"30" => DATA <= x"00";
      when x"31" => DATA <= x"00";
      when x"32" => DATA <= x"00";
      when x"33" => DATA <= x"1C";
      when x"34" => DATA <= x"22";
      when x"35" => DATA <= x"02";
      when x"36" => DATA <= x"04";
      when x"37" => DATA <= x"02";
      when x"38" => DATA <= x"22";
      when x"39" => DATA <= x"1C";
      when x"3A" => DATA <= x"00";
      when x"3B" => DATA <= x"00";
      when x"3C" => DATA <= x"00";
      when x"3D" => DATA <= x"00";
      when x"3E" => DATA <= x"00";
      when x"3F" => DATA <= x"00";
      when x"40" => DATA <= x"00";
      when x"41" => DATA <= x"00";
      when x"42" => DATA <= x"00";
      when x"43" => DATA <= x"04";
      when x"44" => DATA <= x"0C";
      when x"45" => DATA <= x"14";
      when x"46" => DATA <= x"3E";
      when x"47" => DATA <= x"04";
      when x"48" => DATA <= x"04";
      when x"49" => DATA <= x"04";
      when x"4A" => DATA <= x"00";
      when x"4B" => DATA <= x"00";
      when x"4C" => DATA <= x"00";
      when x"4D" => DATA <= x"00";
      when x"4E" => DATA <= x"00";
      when x"4F" => DATA <= x"00";
      when x"50" => DATA <= x"00";
      when x"51" => DATA <= x"00";
      when x"52" => DATA <= x"00";
      when x"53" => DATA <= x"3E";
      when x"54" => DATA <= x"20";
      when x"55" => DATA <= x"3C";
      when x"56" => DATA <= x"02";
      when x"57" => DATA <= x"02";
      when x"58" => DATA <= x"22";
      when x"59" => DATA <= x"1C";
      when x"5A" => DATA <= x"00";
      when x"5B" => DATA <= x"00";
      when x"5C" => DATA <= x"00";
      when x"5D" => DATA <= x"00";
      when x"5E" => DATA <= x"00";
      when x"5F" => DATA <= x"00";
      when x"60" => DATA <= x"00";
      when x"61" => DATA <= x"00";
      when x"62" => DATA <= x"00";
      when x"63" => DATA <= x"1C";
      when x"64" => DATA <= x"20";
      when x"65" => DATA <= x"20";
      when x"66" => DATA <= x"3C";
      when x"67" => DATA <= x"22";
      when x"68" => DATA <= x"22";
      when x"69" => DATA <= x"1C";
      when x"6A" => DATA <= x"00";
      when x"6B" => DATA <= x"00";
      when x"6C" => DATA <= x"00";
      when x"6D" => DATA <= x"00";
      when x"6E" => DATA <= x"00";
      when x"6F" => DATA <= x"00";
      when x"70" => DATA <= x"00";
      when x"71" => DATA <= x"00";
      when x"72" => DATA <= x"00";
      when x"73" => DATA <= x"3E";
      when x"74" => DATA <= x"02";
      when x"75" => DATA <= x"04";
      when x"76" => DATA <= x"08";
      when x"77" => DATA <= x"10";
      when x"78" => DATA <= x"20";
      when x"79" => DATA <= x"20";
      when x"7A" => DATA <= x"00";
      when x"7B" => DATA <= x"00";
      when x"7C" => DATA <= x"00";
      when x"7D" => DATA <= x"00";
      when x"7E" => DATA <= x"00";
      when x"7F" => DATA <= x"00";
      when x"80" => DATA <= x"00";
      when x"81" => DATA <= x"00";
      when x"82" => DATA <= x"00";
      when x"83" => DATA <= x"1C";
      when x"84" => DATA <= x"22";
      when x"85" => DATA <= x"22";
      when x"86" => DATA <= x"1C";
      when x"87" => DATA <= x"22";
      when x"88" => DATA <= x"22";
      when x"89" => DATA <= x"1C";
      when x"8A" => DATA <= x"00";
      when x"8B" => DATA <= x"00";
      when x"8C" => DATA <= x"00";
      when x"8D" => DATA <= x"00";
      when x"8E" => DATA <= x"00";
      when x"8F" => DATA <= x"00";
      when x"90" => DATA <= x"00";
      when x"91" => DATA <= x"00";
      when x"92" => DATA <= x"00";
      when x"93" => DATA <= x"1C";
      when x"94" => DATA <= x"22";
      when x"95" => DATA <= x"22";
      when x"96" => DATA <= x"1E";
      when x"97" => DATA <= x"02";
      when x"98" => DATA <= x"02";
      when x"99" => DATA <= x"1C";
      when x"9A" => DATA <= x"00";
      when x"9B" => DATA <= x"00";
      when x"9C" => DATA <= x"00";
      when x"9D" => DATA <= x"00";
      when x"9E" => DATA <= x"00";
      when x"9F" => DATA <= x"00";
      when x"A0" => DATA <= x"00";
      when x"A1" => DATA <= x"00";
      when x"A2" => DATA <= x"00";
      when x"A3" => DATA <= x"00";
      when x"A4" => DATA <= x"18";
      when x"A5" => DATA <= x"18";
      when x"A6" => DATA <= x"00";
      when x"A7" => DATA <= x"18";
      when x"A8" => DATA <= x"18";
      when x"A9" => DATA <= x"00";
      when x"AA" => DATA <= x"00";
      when x"AB" => DATA <= x"00";
      when x"AC" => DATA <= x"00";
      when x"AD" => DATA <= x"00";
      when x"AE" => DATA <= x"00";
      when x"AF" => DATA <= x"00";
      when x"B0" => DATA <= x"00";
      when x"B1" => DATA <= x"00";
      when x"B2" => DATA <= x"00";
      when x"B3" => DATA <= x"18";
      when x"B4" => DATA <= x"18";
      when x"B5" => DATA <= x"00";
      when x"B6" => DATA <= x"18";
      when x"B7" => DATA <= x"18";
      when x"B8" => DATA <= x"08";
      when x"B9" => DATA <= x"10";
      when x"BA" => DATA <= x"00";
      when x"BB" => DATA <= x"00";
      when x"BC" => DATA <= x"00";
      when x"BD" => DATA <= x"00";
      when x"BE" => DATA <= x"00";
      when x"BF" => DATA <= x"00";
      when x"C0" => DATA <= x"00";
      when x"C1" => DATA <= x"00";
      when x"C2" => DATA <= x"00";
      when x"C3" => DATA <= x"04";
      when x"C4" => DATA <= x"08";
      when x"C5" => DATA <= x"10";
      when x"C6" => DATA <= x"20";
      when x"C7" => DATA <= x"10";
      when x"C8" => DATA <= x"08";
      when x"C9" => DATA <= x"04";
      when x"CA" => DATA <= x"00";
      when x"CB" => DATA <= x"00";
      when x"CC" => DATA <= x"00";
      when x"CD" => DATA <= x"00";
      when x"CE" => DATA <= x"00";
      when x"CF" => DATA <= x"00";
      when x"D0" => DATA <= x"00";
      when x"D1" => DATA <= x"00";
      when x"D2" => DATA <= x"00";
      when x"D3" => DATA <= x"00";
      when x"D4" => DATA <= x"00";
      when x"D5" => DATA <= x"3E";
      when x"D6" => DATA <= x"00";
      when x"D7" => DATA <= x"3E";
      when x"D8" => DATA <= x"00";
      when x"D9" => DATA <= x"00";
      when x"DA" => DATA <= x"00";
      when x"DB" => DATA <= x"00";
      when x"DC" => DATA <= x"00";
      when x"DD" => DATA <= x"00";
      when x"DE" => DATA <= x"00";
      when x"DF" => DATA <= x"00";
      when x"E0" => DATA <= x"00";
      when x"E1" => DATA <= x"00";
      when x"E2" => DATA <= x"00";
      when x"E3" => DATA <= x"10";
      when x"E4" => DATA <= x"08";
      when x"E5" => DATA <= x"04";
      when x"E6" => DATA <= x"02";
      when x"E7" => DATA <= x"04";
      when x"E8" => DATA <= x"08";
      when x"E9" => DATA <= x"10";
      when x"EA" => DATA <= x"00";
      when x"EB" => DATA <= x"00";
      when x"EC" => DATA <= x"00";
      when x"ED" => DATA <= x"00";
      when x"EE" => DATA <= x"00";
      when x"EF" => DATA <= x"00";
      when x"F0" => DATA <= x"00";
      when x"F1" => DATA <= x"00";
      when x"F2" => DATA <= x"00";
      when x"F3" => DATA <= x"18";
      when x"F4" => DATA <= x"24";
      when x"F5" => DATA <= x"04";
      when x"F6" => DATA <= x"08";
      when x"F7" => DATA <= x"08";
      when x"F8" => DATA <= x"00";
      when x"F9" => DATA <= x"08";
      when x"FA" => DATA <= x"00";
      when x"FB" => DATA <= x"00";
      when x"FC" => DATA <= x"00";
      when x"FD" => DATA <= x"00";
      when x"FE" => DATA <= x"00";
      when x"FF" => DATA <= x"00";
      when others => DATA <= (others => '0');
    end case;
	 end if;
  end process;
end RTL;
