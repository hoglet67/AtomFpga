library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- This contains 2.C of the AtoMMC2 firmware (10K x 16)

-- For f_log2 definition
use WORK.SynthCtrlPack.all;

entity XPM is
    generic (
        WIDTH : integer;
        SIZE  : integer
    );
    port(
        cp2     : in  std_logic;
        ce      : in  std_logic;
        address : in  std_logic_vector(f_log2(SIZE) - 1 downto 0);
        din     : in  std_logic_vector(WIDTH - 1 downto 0);
        dout    : out std_logic_vector(WIDTH - 1 downto 0);
        we      : in  std_logic
    );
end;

architecture RTL of XPM is

    type ram_type is array (0 to SIZE - 1) of std_logic_vector (WIDTH - 1 downto 0);

    signal RAM : ram_type := (
        x"940C",
        x"003D",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"009B",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"940C",
        x"005F",
        x"4F42",
        x"544F",
        x"5244",
        x"2E56",
        x"4643",
        x"0047",
        x"4F42",
        x"544F",
        x"5244",
        x"2E56",
        x"4643",
        x"0047",
        x"002A",
        x"2411",
        x"BE1F",
        x"EFCF",
        x"E0DF",
        x"BFDE",
        x"BFCD",
        x"E010",
        x"E6A0",
        x"E0B0",
        x"EBE4",
        x"E4F7",
        x"EF0F",
        x"9503",
        x"BF0B",
        x"C004",
        x"95D8",
        x"920D",
        x"9631",
        x"F3C8",
        x"39AE",
        x"07B1",
        x"F7C9",
        x"E02D",
        x"E9AE",
        x"E0B0",
        x"C001",
        x"921D",
        x"33A6",
        x"07B2",
        x"F7E1",
        x"940E",
        x"2287",
        x"940C",
        x"23D8",
        x"940C",
        x"0000",
        x"E020",
        x"E030",
        x"2E08",
        x"0C00",
        x"0B99",
        x"1728",
        x"0739",
        x"F42C",
        x"98C7",
        x"9AC7",
        x"5F2F",
        x"4F3F",
        x"CFF8",
        x"9508",
        x"E020",
        x"E030",
        x"2E08",
        x"0C00",
        x"0B99",
        x"1728",
        x"0739",
        x"F42C",
        x"98C6",
        x"9AC6",
        x"5F2F",
        x"4F3F",
        x"CFF8",
        x"9508",
        x"2F18",
        x"9AC6",
        x"E1C9",
        x"E0D0",
        x"2F81",
        x"940E",
        x"0061",
        x"9721",
        x"F7D9",
        x"CFFF",
        x"BA1A",
        x"B78A",
        x"7F8C",
        x"BF8A",
        x"B78A",
        x"6082",
        x"BF8A",
        x"B789",
        x"7F8C",
        x"BF89",
        x"98BC",
        x"9AC4",
        x"9AB8",
        x"9AC0",
        x"9AB9",
        x"9AC1",
        x"9ABB",
        x"98C3",
        x"988B",
        x"9508",
        x"921F",
        x"920F",
        x"B60F",
        x"920F",
        x"2411",
        x"900F",
        x"BE0F",
        x"900F",
        x"901F",
        x"9518",
        x"9A8B",
        x"9893",
        x"E98F",
        x"E09F",
        x"9701",
        x"F7F1",
        x"C000",
        x"0000",
        x"988B",
        x"9893",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"0F48",
        x"1F59",
        x"1784",
        x"0795",
        x"F039",
        x"9121",
        x"2FA8",
        x"2FB9",
        x"932D",
        x"2F8A",
        x"2F9B",
        x"CFF6",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2EE6",
        x"2EF7",
        x"E029",
        x"0EE2",
        x"1CF1",
        x"2FA8",
        x"2FB9",
        x"961E",
        x"910D",
        x"911D",
        x"912D",
        x"913C",
        x"9751",
        x"1501",
        x"0511",
        x"0521",
        x"0531",
        x"F409",
        x"C060",
        x"9652",
        x"91CD",
        x"91DC",
        x"9753",
        x"2F2C",
        x"2F3D",
        x"2FE6",
        x"2FF7",
        x"9671",
        x"2FA2",
        x"2FB3",
        x"918D",
        x"2F2A",
        x"2F3B",
        x"3280",
        x"F089",
        x"3085",
        x"F409",
        x"EE85",
        x"EFBF",
        x"1AEB",
        x"0AFB",
        x"2D4E",
        x"2D5F",
        x"5041",
        x"0951",
        x"2FA4",
        x"2FB5",
        x"938C",
        x"16EE",
        x"06FF",
        x"F749",
        x"C002",
        x"2DEE",
        x"2DFF",
        x"8588",
        x"3280",
        x"F0E9",
        x"E28E",
        x"8380",
        x"2F0C",
        x"2F1D",
        x"5F08",
        x"4F1F",
        x"2F2E",
        x"2F3F",
        x"5F2C",
        x"4F3F",
        x"9631",
        x"2FA0",
        x"2FB1",
        x"918D",
        x"2F0A",
        x"2F1B",
        x"3280",
        x"F059",
        x"9631",
        x"2F4E",
        x"2F5F",
        x"5041",
        x"0951",
        x"2FA4",
        x"2FB5",
        x"938C",
        x"17E2",
        x"07F3",
        x"F771",
        x"858B",
        x"2FA6",
        x"2FB7",
        x"9618",
        x"938C",
        x"9718",
        x"8D0C",
        x"8D1D",
        x"8D2E",
        x"8D3F",
        x"930D",
        x"931D",
        x"932D",
        x"933C",
        x"9713",
        x"8D88",
        x"8D99",
        x"9615",
        x"939C",
        x"938E",
        x"9714",
        x"898E",
        x"899F",
        x"9617",
        x"939C",
        x"938E",
        x"9716",
        x"2EEE",
        x"2EFF",
        x"2DEE",
        x"2DFF",
        x"8210",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"2331",
        x"E0A0",
        x"E0B0",
        x"E5E2",
        x"E0F1",
        x"940C",
        x"230F",
        x"2FE8",
        x"2FF9",
        x"A486",
        x"A497",
        x"A8A0",
        x"A8B1",
        x"1684",
        x"0695",
        x"06A6",
        x"06B7",
        x"F409",
        x"C058",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"2FC8",
        x"2FD9",
        x"8184",
        x"2388",
        x"F439",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F409",
        x"C049",
        x"C038",
        x"A962",
        x"A973",
        x"E001",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"8181",
        x"940E",
        x"1846",
        x"2B89",
        x"F019",
        x"E081",
        x"E090",
        x"C03B",
        x"821C",
        x"8D4A",
        x"8D5B",
        x"8D6C",
        x"8D7D",
        x"A18A",
        x"A19B",
        x"A1AC",
        x"A1BD",
        x"0F84",
        x"1F95",
        x"1FA6",
        x"1FB7",
        x"1688",
        x"0699",
        x"06AA",
        x"06BB",
        x"F6C0",
        x"811B",
        x"3012",
        x"F2A8",
        x"8D8A",
        x"8D9B",
        x"8DAC",
        x"8DBD",
        x"0E88",
        x"1E99",
        x"1EAA",
        x"1EBB",
        x"A96A",
        x"A97B",
        x"E001",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"8189",
        x"940E",
        x"1846",
        x"5011",
        x"CFEA",
        x"A96A",
        x"A97B",
        x"E001",
        x"2D5F",
        x"2D4E",
        x"2D3D",
        x"2D2C",
        x"8189",
        x"940E",
        x"183C",
        x"2B89",
        x"F641",
        x"A6CE",
        x"A6DF",
        x"AAE8",
        x"AAF9",
        x"E080",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"232B",
        x"930F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F24",
        x"2F35",
        x"2F46",
        x"2F57",
        x"A96A",
        x"A97B",
        x"E001",
        x"8189",
        x"940E",
        x"183C",
        x"2B89",
        x"F519",
        x"A9EA",
        x"A9FB",
        x"2FAE",
        x"2FBF",
        x"50A2",
        x"4FBE",
        x"918D",
        x"919C",
        x"3585",
        x"4A9A",
        x"F4D1",
        x"A986",
        x"A997",
        x"ADA0",
        x"ADB1",
        x"27BB",
        x"3486",
        x"4491",
        x"45A4",
        x"05B1",
        x"F091",
        x"5AEE",
        x"4FFF",
        x"8140",
        x"8151",
        x"8162",
        x"8173",
        x"2777",
        x"E081",
        x"3446",
        x"4451",
        x"4564",
        x"0571",
        x"F431",
        x"C004",
        x"E083",
        x"C003",
        x"E082",
        x"C001",
        x"E080",
        x"91DF",
        x"91CF",
        x"910F",
        x"9508",
        x"9700",
        x"F091",
        x"2FE8",
        x"2FF9",
        x"8120",
        x"2322",
        x"F069",
        x"8126",
        x"8137",
        x"1726",
        x"0737",
        x"F441",
        x"8181",
        x"940E",
        x"1839",
        x"FD80",
        x"C006",
        x"E080",
        x"E090",
        x"9508",
        x"E089",
        x"E090",
        x"9508",
        x"E083",
        x"E090",
        x"9508",
        x"930F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"940E",
        x"014C",
        x"9700",
        x"F009",
        x"C05C",
        x"8188",
        x"3083",
        x"F009",
        x"C04B",
        x"818D",
        x"2388",
        x"F409",
        x"C047",
        x"A61E",
        x"A61F",
        x"AA18",
        x"AA19",
        x"A9EA",
        x"A9FB",
        x"2F8E",
        x"2F9F",
        x"5F9E",
        x"17E8",
        x"07F9",
        x"F011",
        x"9211",
        x"CFFB",
        x"A96A",
        x"A97B",
        x"2FE6",
        x"2FF7",
        x"50E2",
        x"4FFE",
        x"E585",
        x"EA9A",
        x"8391",
        x"8380",
        x"E582",
        x"E592",
        x"E6A1",
        x"E4B1",
        x"2FE6",
        x"2FF7",
        x"8380",
        x"8391",
        x"83A2",
        x"83B3",
        x"51EC",
        x"4FFE",
        x"E782",
        x"E792",
        x"E4A1",
        x"E6B1",
        x"8380",
        x"8391",
        x"83A2",
        x"83B3",
        x"858E",
        x"859F",
        x"89A8",
        x"89B9",
        x"9634",
        x"8380",
        x"8391",
        x"83A2",
        x"83B3",
        x"858A",
        x"859B",
        x"85AC",
        x"85BD",
        x"9634",
        x"8380",
        x"8391",
        x"83A2",
        x"83B3",
        x"892A",
        x"893B",
        x"894C",
        x"895D",
        x"E001",
        x"8189",
        x"940E",
        x"1846",
        x"821D",
        x"E040",
        x"E050",
        x"E060",
        x"8189",
        x"940E",
        x"1850",
        x"E031",
        x"E020",
        x"2B89",
        x"F409",
        x"E030",
        x"2F83",
        x"2F92",
        x"91DF",
        x"91CF",
        x"910F",
        x"9508",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"C0A9",
        x"8D8E",
        x"8D9F",
        x"A1A8",
        x"A1B9",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C09F",
        x"A04A",
        x"A05B",
        x"A06C",
        x"A07D",
        x"8188",
        x"3082",
        x"F409",
        x"C053",
        x"3083",
        x"F409",
        x"C06D",
        x"3081",
        x"F009",
        x"C096",
        x"2EA4",
        x"2EB5",
        x"94B6",
        x"94A7",
        x"0CAC",
        x"1CBD",
        x"2D8A",
        x"2D9B",
        x"2F89",
        x"2799",
        x"9586",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"014C",
        x"2B89",
        x"F009",
        x"C07C",
        x"2D8A",
        x"2D9B",
        x"7091",
        x"A9EA",
        x"A9FB",
        x"0FE8",
        x"1FF9",
        x"8110",
        x"EF8F",
        x"1AA8",
        x"0AB8",
        x"2D8A",
        x"2D9B",
        x"2F89",
        x"2799",
        x"9586",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"014C",
        x"2B89",
        x"F009",
        x"C05D",
        x"E081",
        x"22B8",
        x"A9EA",
        x"A9FB",
        x"0DEA",
        x"1DFB",
        x"8180",
        x"2F61",
        x"E070",
        x"2B78",
        x"FEC0",
        x"C006",
        x"E044",
        x"9576",
        x"9567",
        x"954A",
        x"F7E1",
        x"C01C",
        x"707F",
        x"C01A",
        x"2F45",
        x"2F56",
        x"2F67",
        x"2777",
        x"0D44",
        x"1D55",
        x"1D66",
        x"1D77",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"014C",
        x"2B89",
        x"F5D9",
        x"0CCC",
        x"1CDD",
        x"94E8",
        x"F8C0",
        x"E081",
        x"22D8",
        x"A9EA",
        x"A9FB",
        x"0DEC",
        x"1DFD",
        x"8160",
        x"8171",
        x"E080",
        x"E090",
        x"C030",
        x"E097",
        x"9576",
        x"9567",
        x"9557",
        x"9547",
        x"959A",
        x"F7D1",
        x"0D44",
        x"1D55",
        x"1D66",
        x"1D77",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"014C",
        x"2B89",
        x"F4D9",
        x"0CCC",
        x"1CDD",
        x"0CCC",
        x"1CDD",
        x"EF8C",
        x"22C8",
        x"E081",
        x"22D8",
        x"A9EA",
        x"A9FB",
        x"0DEC",
        x"1DFD",
        x"8180",
        x"8191",
        x"81A2",
        x"81B3",
        x"2F68",
        x"2F79",
        x"2F8A",
        x"2F9B",
        x"709F",
        x"C009",
        x"E061",
        x"E070",
        x"E080",
        x"E090",
        x"C004",
        x"EF6F",
        x"EF7F",
        x"EF8F",
        x"EF9F",
        x"91DF",
        x"91CF",
        x"911F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"9508",
        x"E0A8",
        x"E0B0",
        x"E6E1",
        x"E0F3",
        x"940C",
        x"230B",
        x"2E88",
        x"2E99",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"8309",
        x"831A",
        x"832B",
        x"833C",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"C0F2",
        x"2FE8",
        x"2FF9",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C0E6",
        x"A042",
        x"A053",
        x"A064",
        x"A075",
        x"8180",
        x"3082",
        x"F409",
        x"C08A",
        x"3083",
        x"F409",
        x"C0A9",
        x"3081",
        x"F009",
        x"C0D0",
        x"2EA4",
        x"2EB5",
        x"94B6",
        x"94A7",
        x"0EA4",
        x"1EB5",
        x"2D8A",
        x"2D9B",
        x"2F89",
        x"2799",
        x"9586",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2D88",
        x"2D99",
        x"940E",
        x"014C",
        x"9700",
        x"F009",
        x"C0B8",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"2D8A",
        x"2D9B",
        x"7091",
        x"2F2E",
        x"2F3F",
        x"0F28",
        x"1F39",
        x"2DBF",
        x"2DAE",
        x"2D9D",
        x"2D8C",
        x"7081",
        x"2799",
        x"27AA",
        x"27BB",
        x"838D",
        x"839E",
        x"83AF",
        x"87B8",
        x"FEC0",
        x"C009",
        x"2FA2",
        x"2FB3",
        x"918C",
        x"708F",
        x"8199",
        x"9592",
        x"7F90",
        x"2B89",
        x"C001",
        x"8189",
        x"2FE2",
        x"2FF3",
        x"8380",
        x"EFFF",
        x"1AAF",
        x"0ABF",
        x"E081",
        x"2DA8",
        x"2DB9",
        x"9614",
        x"938C",
        x"2D8A",
        x"2D9B",
        x"2F89",
        x"2799",
        x"9586",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"0F48",
        x"1F59",
        x"1D61",
        x"1D71",
        x"2D88",
        x"2D99",
        x"940E",
        x"014C",
        x"9700",
        x"F009",
        x"C074",
        x"E0B1",
        x"22BB",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"0DEA",
        x"1DFB",
        x"812D",
        x"813E",
        x"814F",
        x"8558",
        x"2B23",
        x"2B24",
        x"2B25",
        x"F061",
        x"8049",
        x"805A",
        x"806B",
        x"807C",
        x"E064",
        x"9476",
        x"9467",
        x"9457",
        x"9447",
        x"956A",
        x"F7D1",
        x"C006",
        x"8130",
        x"7F30",
        x"812A",
        x"702F",
        x"2E43",
        x"2A42",
        x"8240",
        x"C04E",
        x"2777",
        x"2D6F",
        x"2D5E",
        x"2D4D",
        x"0D44",
        x"1D55",
        x"1D66",
        x"1D77",
        x"2D88",
        x"2D99",
        x"940E",
        x"014C",
        x"9700",
        x"F009",
        x"C03F",
        x"0CCC",
        x"1CDD",
        x"94E8",
        x"F8C0",
        x"E031",
        x"22D3",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"0DEC",
        x"1DFD",
        x"8129",
        x"813A",
        x"8331",
        x"8320",
        x"C02C",
        x"E037",
        x"9576",
        x"9567",
        x"9557",
        x"9547",
        x"953A",
        x"F7D1",
        x"0D44",
        x"1D55",
        x"1D66",
        x"1D77",
        x"2D88",
        x"2D99",
        x"940E",
        x"014C",
        x"9700",
        x"F4D9",
        x"0CCC",
        x"1CDD",
        x"0CCC",
        x"1CDD",
        x"EF3C",
        x"22C3",
        x"E031",
        x"22D3",
        x"2DA8",
        x"2DB9",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"0DEC",
        x"1DFD",
        x"8129",
        x"813A",
        x"814B",
        x"815C",
        x"8320",
        x"8331",
        x"8342",
        x"8353",
        x"C002",
        x"E082",
        x"E090",
        x"E021",
        x"2DA8",
        x"2DB9",
        x"9614",
        x"932C",
        x"C002",
        x"E082",
        x"E090",
        x"9628",
        x"E1E0",
        x"940C",
        x"2327",
        x"E0A4",
        x"E0B0",
        x"E6EF",
        x"E0F4",
        x"940C",
        x"2309",
        x"2E28",
        x"2E39",
        x"2E44",
        x"2E55",
        x"2E66",
        x"2E77",
        x"2FA8",
        x"2FB9",
        x"965E",
        x"912D",
        x"913D",
        x"914D",
        x"915C",
        x"9791",
        x"8329",
        x"833A",
        x"834B",
        x"835C",
        x"1441",
        x"0451",
        x"0461",
        x"0471",
        x"F489",
        x"961A",
        x"908D",
        x"909D",
        x"90AD",
        x"90BC",
        x"971D",
        x"1481",
        x"0491",
        x"04A1",
        x"04B1",
        x"F109",
        x"1682",
        x"0693",
        x"06A4",
        x"06B5",
        x"F108",
        x"C01B",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"940E",
        x"0282",
        x"3062",
        x"0571",
        x"0581",
        x"0591",
        x"F408",
        x"C09F",
        x"8129",
        x"813A",
        x"814B",
        x"815C",
        x"1762",
        x"0773",
        x"0784",
        x"0795",
        x"F408",
        x"C09A",
        x"2CB7",
        x"2CA6",
        x"2C95",
        x"2C84",
        x"C005",
        x"2488",
        x"9483",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"2CFB",
        x"2CEA",
        x"2CD9",
        x"2CC8",
        x"EF3F",
        x"1AC3",
        x"0AD3",
        x"0AE3",
        x"0AF3",
        x"8129",
        x"813A",
        x"814B",
        x"815C",
        x"16C2",
        x"06D3",
        x"06E4",
        x"06F5",
        x"F068",
        x"E032",
        x"1683",
        x"0491",
        x"04A1",
        x"04B1",
        x"F410",
        x"E040",
        x"C072",
        x"E082",
        x"2EC8",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2D82",
        x"2D93",
        x"940E",
        x"0282",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F099",
        x"3F6F",
        x"EF4F",
        x"0774",
        x"0784",
        x"0794",
        x"F409",
        x"C05D",
        x"3061",
        x"0571",
        x"0581",
        x"0591",
        x"F409",
        x"C057",
        x"14C8",
        x"04D9",
        x"04EA",
        x"04FB",
        x"F631",
        x"CFD9",
        x"EF0F",
        x"EF1F",
        x"EF2F",
        x"E03F",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2D82",
        x"2D93",
        x"940E",
        x"035B",
        x"2B89",
        x"F029",
        x"EF4F",
        x"EF3F",
        x"EF2F",
        x"EF9F",
        x"C041",
        x"1441",
        x"0451",
        x"0461",
        x"0471",
        x"F501",
        x"2DA2",
        x"2DB3",
        x"961A",
        x"92CD",
        x"92DD",
        x"92ED",
        x"92FC",
        x"971D",
        x"961E",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"3F8F",
        x"EFEF",
        x"079E",
        x"07AE",
        x"07BE",
        x"F0D9",
        x"9701",
        x"09A1",
        x"09B1",
        x"2DE2",
        x"2DF3",
        x"8786",
        x"8797",
        x"8BA0",
        x"8BB1",
        x"E081",
        x"8385",
        x"C00F",
        x"2D3F",
        x"2D2E",
        x"2D1D",
        x"2D0C",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"2D82",
        x"2D93",
        x"940E",
        x"035B",
        x"2B89",
        x"F641",
        x"CFD1",
        x"2D4C",
        x"2D3D",
        x"2D2E",
        x"2D9F",
        x"C008",
        x"E041",
        x"E030",
        x"E020",
        x"E090",
        x"C003",
        x"2F46",
        x"2F37",
        x"2F28",
        x"2F64",
        x"2F73",
        x"2F82",
        x"9624",
        x"E1E2",
        x"940C",
        x"2325",
        x"E0A0",
        x"E0B0",
        x"E5E7",
        x"E0F5",
        x"940C",
        x"230E",
        x"2FC8",
        x"2FD9",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F418",
        x"E082",
        x"E090",
        x"C05A",
        x"8D8E",
        x"8D9F",
        x"A1A8",
        x"A1B9",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F7A0",
        x"2477",
        x"9473",
        x"8D8E",
        x"8D9F",
        x"A1A8",
        x"A1B9",
        x"16C8",
        x"06D9",
        x"06EA",
        x"06FB",
        x"F480",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"0282",
        x"2E86",
        x"2E97",
        x"2EA8",
        x"2EB9",
        x"2B67",
        x"2B68",
        x"2B69",
        x"F419",
        x"E080",
        x"E090",
        x"C033",
        x"E081",
        x"1688",
        x"0491",
        x"04A1",
        x"04B1",
        x"F281",
        x"EF2F",
        x"1682",
        x"0692",
        x"06A2",
        x"06B2",
        x"F129",
        x"E000",
        x"E010",
        x"E020",
        x"E030",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"035B",
        x"9700",
        x"F4C9",
        x"858E",
        x"859F",
        x"89A8",
        x"89B9",
        x"3F8F",
        x"EF2F",
        x"0792",
        x"07A2",
        x"07B2",
        x"F041",
        x"9601",
        x"1DA1",
        x"1DB1",
        x"878E",
        x"879F",
        x"8BA8",
        x"8BB9",
        x"827D",
        x"2CFB",
        x"2CEA",
        x"2CD9",
        x"2CC8",
        x"CFB3",
        x"E081",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0ED",
        x"940C",
        x"232A",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F97",
        x"2F86",
        x"2F75",
        x"2F64",
        x"5062",
        x"0971",
        x"0981",
        x"0991",
        x"8CCE",
        x"8CDF",
        x"A0E8",
        x"A0F9",
        x"E022",
        x"1AC2",
        x"08D1",
        x"08E1",
        x"08F1",
        x"156C",
        x"057D",
        x"058E",
        x"059F",
        x"F4B8",
        x"812A",
        x"E030",
        x"E040",
        x"E050",
        x"940E",
        x"22E5",
        x"2E82",
        x"2E93",
        x"2EA4",
        x"2EB5",
        x"A58A",
        x"A59B",
        x"A5AC",
        x"A5BD",
        x"2F68",
        x"2F79",
        x"2F8A",
        x"2F9B",
        x"0D68",
        x"1D79",
        x"1D8A",
        x"1D9B",
        x"C004",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2FC6",
        x"2FD7",
        x"2FA8",
        x"2FB9",
        x"9615",
        x"937C",
        x"936E",
        x"9714",
        x"9616",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9719",
        x"3041",
        x"0551",
        x"0561",
        x"0571",
        x"F419",
        x"E082",
        x"E090",
        x"C09D",
        x"2FA8",
        x"2FB9",
        x"91ED",
        x"91FC",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F780",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F529",
        x"8180",
        x"3083",
        x"F449",
        x"A146",
        x"A157",
        x"A560",
        x"A571",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F4C9",
        x"2FA0",
        x"2FB1",
        x"961A",
        x"921D",
        x"921D",
        x"921D",
        x"921C",
        x"971D",
        x"8580",
        x"8591",
        x"17C8",
        x"07D9",
        x"F690",
        x"A186",
        x"A197",
        x"A5A0",
        x"A5B1",
        x"2F2C",
        x"2F3D",
        x"E0F4",
        x"9536",
        x"9527",
        x"95FA",
        x"F7E1",
        x"C043",
        x"80E2",
        x"2CF1",
        x"E0E4",
        x"0CEE",
        x"1CFF",
        x"95EA",
        x"F7E1",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"8191",
        x"15CE",
        x"05DF",
        x"F120",
        x"940E",
        x"0282",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"3F4F",
        x"EFFF",
        x"075F",
        x"076F",
        x"077F",
        x"F409",
        x"C049",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"CFA5",
        x"2FA0",
        x"2FB1",
        x"91ED",
        x"91FC",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"CF97",
        x"19CE",
        x"09DF",
        x"CFD5",
        x"8742",
        x"8753",
        x"8764",
        x"8775",
        x"940E",
        x"05C4",
        x"2F2C",
        x"2F3D",
        x"E044",
        x"9536",
        x"9527",
        x"954A",
        x"F7E1",
        x"2FB9",
        x"2FA8",
        x"2F97",
        x"2F86",
        x"0F82",
        x"1F93",
        x"1DA1",
        x"1DB1",
        x"2FE0",
        x"2FF1",
        x"8786",
        x"8797",
        x"8BA0",
        x"8BB1",
        x"2FA0",
        x"2FB1",
        x"9001",
        x"81F0",
        x"2DE0",
        x"70CF",
        x"27DD",
        x"E085",
        x"0FCC",
        x"1FDD",
        x"958A",
        x"F7E1",
        x"A982",
        x"A993",
        x"0FC8",
        x"1FD9",
        x"9653",
        x"93DC",
        x"93CE",
        x"9752",
        x"E080",
        x"E090",
        x"C002",
        x"E081",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"2331",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"816C",
        x"817D",
        x"940E",
        x"060C",
        x"9700",
        x"F491",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"9700",
        x"F441",
        x"89EA",
        x"89FB",
        x"EE25",
        x"8320",
        x"81E8",
        x"81F9",
        x"E021",
        x"8324",
        x"91DF",
        x"91CF",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"EFE1",
        x"E0F6",
        x"940C",
        x"230F",
        x"2FC8",
        x"2FD9",
        x"2EC6",
        x"2ED7",
        x"810C",
        x"811D",
        x"5F0F",
        x"4F1F",
        x"F419",
        x"E084",
        x"E090",
        x"C0FB",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F3A1",
        x"2EE0",
        x"2EF1",
        x"E08F",
        x"22E8",
        x"24FF",
        x"14E1",
        x"04F1",
        x"F009",
        x"C0D5",
        x"5F4F",
        x"4F5F",
        x"4F6F",
        x"4F7F",
        x"874E",
        x"875F",
        x"8B68",
        x"8B79",
        x"854A",
        x"855B",
        x"856C",
        x"857D",
        x"8188",
        x"8199",
        x"2FE8",
        x"2FF9",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F431",
        x"8580",
        x"8591",
        x"1708",
        x"0719",
        x"F688",
        x"C0BA",
        x"8122",
        x"E030",
        x"5021",
        x"0931",
        x"2FE0",
        x"2FF1",
        x"E0A4",
        x"95F6",
        x"95E7",
        x"95AA",
        x"F7E1",
        x"232E",
        x"233F",
        x"2B23",
        x"F009",
        x"C0AA",
        x"940E",
        x"0282",
        x"2E86",
        x"2E97",
        x"2EA8",
        x"2EB9",
        x"3062",
        x"0571",
        x"0581",
        x"0591",
        x"F418",
        x"E082",
        x"E090",
        x"C0B0",
        x"EF8F",
        x"1688",
        x"0698",
        x"06A8",
        x"06B8",
        x"F419",
        x"E081",
        x"E090",
        x"C0A7",
        x"8188",
        x"8199",
        x"2FE8",
        x"2FF9",
        x"8D46",
        x"8D57",
        x"A160",
        x"A171",
        x"1684",
        x"0695",
        x"06A6",
        x"06B7",
        x"F408",
        x"C075",
        x"14C1",
        x"04D1",
        x"F409",
        x"CF97",
        x"854A",
        x"855B",
        x"856C",
        x"857D",
        x"940E",
        x"0469",
        x"2E86",
        x"2E97",
        x"2EA8",
        x"2EB9",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F409",
        x"C083",
        x"3061",
        x"0571",
        x"0581",
        x"0591",
        x"F269",
        x"EF8F",
        x"1688",
        x"0698",
        x"06A8",
        x"06B8",
        x"F281",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"2B89",
        x"F631",
        x"81E8",
        x"81F9",
        x"A802",
        x"A9F3",
        x"2DE0",
        x"2F8E",
        x"2F9F",
        x"5F9E",
        x"17E8",
        x"07F9",
        x"F011",
        x"9211",
        x"CFFB",
        x"80C8",
        x"80D9",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"05C4",
        x"2DEC",
        x"2DFD",
        x"A766",
        x"A777",
        x"AB80",
        x"AB91",
        x"2CD1",
        x"24CC",
        x"94C3",
        x"81E8",
        x"81F9",
        x"8182",
        x"16D8",
        x"F4D8",
        x"82C4",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"2B89",
        x"F009",
        x"CF95",
        x"81E8",
        x"81F9",
        x"A586",
        x"A597",
        x"A9A0",
        x"A9B1",
        x"9601",
        x"1DA1",
        x"1DB1",
        x"A786",
        x"A797",
        x"ABA0",
        x"ABB1",
        x"94D3",
        x"CFE0",
        x"A586",
        x"A597",
        x"A9A0",
        x"A9B1",
        x"198D",
        x"0991",
        x"09A1",
        x"09B1",
        x"A786",
        x"A797",
        x"ABA0",
        x"ABB1",
        x"868A",
        x"869B",
        x"86AC",
        x"86BD",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"8188",
        x"8199",
        x"940E",
        x"05C4",
        x"876E",
        x"877F",
        x"8B88",
        x"8B99",
        x"831D",
        x"830C",
        x"81E8",
        x"81F9",
        x"E085",
        x"0CEE",
        x"1CFF",
        x"958A",
        x"F7E1",
        x"A982",
        x"A993",
        x"0EE8",
        x"1EF9",
        x"8AFB",
        x"8AEA",
        x"E080",
        x"E090",
        x"C002",
        x"E087",
        x"E090",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"232B",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"927F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F26",
        x"2F37",
        x"2FA6",
        x"2FB7",
        x"918D",
        x"2F6A",
        x"2F7B",
        x"3280",
        x"F3B9",
        x"2F02",
        x"2F13",
        x"328F",
        x"F011",
        x"358C",
        x"F449",
        x"2F02",
        x"2F13",
        x"5F0F",
        x"4F1F",
        x"821E",
        x"821F",
        x"8618",
        x"8619",
        x"C00A",
        x"81E8",
        x"81F9",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"838E",
        x"839F",
        x"87A8",
        x"87B9",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"3280",
        x"F028",
        x"E2B0",
        x"2EAB",
        x"E085",
        x"2EB8",
        x"C05C",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"060C",
        x"8A1B",
        x"8A1A",
        x"C11E",
        x"89EA",
        x"89FB",
        x"8180",
        x"2388",
        x"F409",
        x"C0E6",
        x"8583",
        x"FD83",
        x"C015",
        x"89AC",
        x"89BD",
        x"2F4E",
        x"2F5F",
        x"5F45",
        x"4F5F",
        x"17E4",
        x"07F5",
        x"F409",
        x"C0DC",
        x"9181",
        x"912D",
        x"2E08",
        x"0C00",
        x"0B99",
        x"1B82",
        x"0991",
        x"FD27",
        x"9593",
        x"2B89",
        x"F389",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"06EB",
        x"9700",
        x"F451",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"9700",
        x"F281",
        x"89EC",
        x"89FD",
        x"8523",
        x"7024",
        x"9700",
        x"F009",
        x"C0BB",
        x"2322",
        x"F009",
        x"C0BE",
        x"89EA",
        x"89FB",
        x"8583",
        x"FF84",
        x"C0BC",
        x"8984",
        x"8995",
        x"E0A0",
        x"E0B0",
        x"2FA8",
        x"2FB9",
        x"2799",
        x"2788",
        x"8D42",
        x"8D53",
        x"E060",
        x"E070",
        x"2B84",
        x"2B95",
        x"2BA6",
        x"2BB7",
        x"838E",
        x"839F",
        x"87A8",
        x"87B9",
        x"89EC",
        x"89FD",
        x"2F4E",
        x"2F5F",
        x"2F8E",
        x"2F9F",
        x"960B",
        x"2FAE",
        x"2FBF",
        x"17A8",
        x"07B9",
        x"F011",
        x"92AD",
        x"CFFB",
        x"2FA0",
        x"2FB1",
        x"918C",
        x"328E",
        x"F051",
        x"2E20",
        x"2E31",
        x"E080",
        x"E090",
        x"E060",
        x"E070",
        x"E028",
        x"E030",
        x"2C91",
        x"C037",
        x"2F60",
        x"2F71",
        x"E020",
        x"E030",
        x"5F2F",
        x"4F3F",
        x"2FA6",
        x"2FB7",
        x"918D",
        x"2F6A",
        x"2F7B",
        x"328E",
        x"F451",
        x"3023",
        x"0531",
        x"F409",
        x"C07D",
        x"2FA4",
        x"2FB5",
        x"938D",
        x"2F4A",
        x"2F5B",
        x"CFED",
        x"328F",
        x"F029",
        x"358C",
        x"F019",
        x"3281",
        x"F008",
        x"C070",
        x"0F02",
        x"1F13",
        x"3281",
        x"F010",
        x"E280",
        x"C001",
        x"E284",
        x"8783",
        x"C04E",
        x"325F",
        x"F199",
        x"355C",
        x"F189",
        x"325E",
        x"F4A9",
        x"3028",
        x"0531",
        x"F009",
        x"C05D",
        x"0C99",
        x"0C99",
        x"E088",
        x"E090",
        x"E02B",
        x"E030",
        x"5F6F",
        x"4F7F",
        x"2DA2",
        x"2DB3",
        x"915D",
        x"2E2A",
        x"2E3B",
        x"2E75",
        x"3251",
        x"F730",
        x"C06A",
        x"1782",
        x"0793",
        x"F00C",
        x"C048",
        x"FD57",
        x"C046",
        x"2EC5",
        x"2CD1",
        x"E9A3",
        x"2EEA",
        x"E0A0",
        x"2EFA",
        x"2DAE",
        x"2DBF",
        x"914D",
        x"2EEA",
        x"2EFB",
        x"2344",
        x"F1E1",
        x"2E44",
        x"0F44",
        x"0855",
        x"144C",
        x"045D",
        x"F799",
        x"C032",
        x"E040",
        x"2B89",
        x"F179",
        x"8180",
        x"3E85",
        x"F409",
        x"82B0",
        x"3028",
        x"0531",
        x"F411",
        x"0C99",
        x"0C99",
        x"2D89",
        x"7083",
        x"3081",
        x"F409",
        x"6140",
        x"2D89",
        x"708C",
        x"3084",
        x"F409",
        x"6048",
        x"0F06",
        x"1F17",
        x"8743",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"060C",
        x"CF38",
        x"E084",
        x"E090",
        x"CF41",
        x"E080",
        x"E090",
        x"CF3E",
        x"3084",
        x"0591",
        x"F549",
        x"2322",
        x"F021",
        x"C026",
        x"E080",
        x"E090",
        x"C023",
        x"E085",
        x"E090",
        x"C020",
        x"E086",
        x"E090",
        x"C01D",
        x"EB4F",
        x"0F45",
        x"314A",
        x"F420",
        x"2DB9",
        x"60B2",
        x"2E9B",
        x"C00A",
        x"E94F",
        x"0F45",
        x"314A",
        x"F430",
        x"2D49",
        x"6041",
        x"2E94",
        x"EE40",
        x"2E74",
        x"0E75",
        x"2F4E",
        x"2F5F",
        x"0F48",
        x"1F59",
        x"2FA4",
        x"2FB5",
        x"927C",
        x"9601",
        x"CF8B",
        x"E044",
        x"CFAF",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"907F",
        x"905F",
        x"904F",
        x"903F",
        x"902F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"E060",
        x"E070",
        x"940E",
        x"060C",
        x"2F08",
        x"2F19",
        x"2B89",
        x"F009",
        x"C045",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"2F08",
        x"2F19",
        x"2B89",
        x"F5C9",
        x"89EA",
        x"89FB",
        x"8180",
        x"3E85",
        x"F049",
        x"2388",
        x"F039",
        x"E061",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"06EB",
        x"CFE1",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"2F08",
        x"2F19",
        x"2B89",
        x"F4F9",
        x"88EA",
        x"88FB",
        x"2DEE",
        x"2DFF",
        x"2D8E",
        x"2D9F",
        x"9680",
        x"17E8",
        x"07F9",
        x"F011",
        x"9211",
        x"CFFB",
        x"896C",
        x"897D",
        x"E04B",
        x"E050",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"00BC",
        x"89EC",
        x"89FD",
        x"8583",
        x"7188",
        x"2DEE",
        x"2DFF",
        x"8784",
        x"81E8",
        x"81F9",
        x"E081",
        x"8384",
        x"2F80",
        x"2F91",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"2331",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"E084",
        x"E090",
        x"854E",
        x"855F",
        x"8968",
        x"8979",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F0E1",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"9700",
        x"F4C1",
        x"89EA",
        x"89FB",
        x"8180",
        x"2388",
        x"F0C1",
        x"3E85",
        x"F031",
        x"8583",
        x"FD83",
        x"C003",
        x"E080",
        x"E090",
        x"C013",
        x"E060",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"06EB",
        x"9700",
        x"F2E1",
        x"C002",
        x"9700",
        x"F391",
        x"861E",
        x"861F",
        x"8A18",
        x"8A19",
        x"C003",
        x"E084",
        x"E090",
        x"CFF8",
        x"91DF",
        x"91CF",
        x"9508",
        x"2F68",
        x"2F79",
        x"EA88",
        x"E093",
        x"940E",
        x"00CB",
        x"9508",
        x"E0A8",
        x"E0B0",
        x"E1E5",
        x"E0FA",
        x"940C",
        x"230A",
        x"2FA8",
        x"2FB9",
        x"91ED",
        x"91FC",
        x"9711",
        x"8120",
        x"2E02",
        x"0C00",
        x"0B33",
        x"5320",
        x"0931",
        x"302A",
        x"0531",
        x"F438",
        x"8151",
        x"335A",
        x"F421",
        x"9632",
        x"93ED",
        x"93FC",
        x"C003",
        x"9120",
        x"009E",
        x"E030",
        x"2B23",
        x"F009",
        x"C1C2",
        x"90C0",
        x"00A1",
        x"90D0",
        x"00A2",
        x"2FE6",
        x"2FF7",
        x"82D1",
        x"82C0",
        x"14C1",
        x"04D1",
        x"F409",
        x"C1B9",
        x"2F14",
        x"2DAC",
        x"2DBD",
        x"918C",
        x"2388",
        x"F071",
        x"9611",
        x"918C",
        x"940E",
        x"1839",
        x"FD80",
        x"C008",
        x"2311",
        x"F409",
        x"C1AD",
        x"FF82",
        x"C1AB",
        x"E08A",
        x"E090",
        x"C1BF",
        x"2DEC",
        x"2DFD",
        x"8210",
        x"8211",
        x"E080",
        x"940E",
        x"1836",
        x"FD80",
        x"C1A2",
        x"2311",
        x"F011",
        x"FD82",
        x"CFF0",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"01BD",
        x"3081",
        x"F509",
        x"2DAC",
        x"2DBD",
        x"96D2",
        x"918D",
        x"919C",
        x"97D3",
        x"2FE8",
        x"2FF9",
        x"53EE",
        x"4FFE",
        x"8120",
        x"2322",
        x"F419",
        x"E08D",
        x"E090",
        x"C198",
        x"2FE8",
        x"2FF9",
        x"53EA",
        x"4FFE",
        x"8080",
        x"8091",
        x"80A2",
        x"80B3",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"01BD",
        x"C004",
        x"2C81",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"3083",
        x"F409",
        x"C16F",
        x"2388",
        x"F719",
        x"2DEC",
        x"2DFD",
        x"A8E2",
        x"A8F3",
        x"2DAE",
        x"2DBF",
        x"961B",
        x"918D",
        x"919C",
        x"971C",
        x"1581",
        x"4092",
        x"F6B1",
        x"2DEE",
        x"2DFF",
        x"8966",
        x"8977",
        x"E080",
        x"E090",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F421",
        x"A164",
        x"A175",
        x"A186",
        x"A197",
        x"2DAC",
        x"2DBD",
        x"965A",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"975D",
        x"2DEE",
        x"2DFF",
        x"8920",
        x"9613",
        x"932C",
        x"E030",
        x"E040",
        x"E050",
        x"940E",
        x"22E5",
        x"8329",
        x"833A",
        x"834B",
        x"835C",
        x"2DAE",
        x"2DBF",
        x"961E",
        x"918D",
        x"919C",
        x"971F",
        x"2C48",
        x"2C59",
        x"2C6A",
        x"2C7B",
        x"0E48",
        x"1E59",
        x"1C61",
        x"1C71",
        x"2DEC",
        x"2DFD",
        x"A242",
        x"A253",
        x"A264",
        x"A275",
        x"961D",
        x"903C",
        x"971D",
        x"8232",
        x"9651",
        x"918D",
        x"919C",
        x"9752",
        x"8791",
        x"8780",
        x"9653",
        x"914D",
        x"915C",
        x"9754",
        x"E060",
        x"E070",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F431",
        x"9690",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9793",
        x"E024",
        x"9596",
        x"9587",
        x"952A",
        x"F7E1",
        x"2F08",
        x"2F19",
        x"E020",
        x"E030",
        x"830D",
        x"831E",
        x"832F",
        x"8738",
        x"2DAE",
        x"2DBF",
        x"961E",
        x"918D",
        x"919C",
        x"971F",
        x"2F04",
        x"2F15",
        x"2F26",
        x"2F37",
        x"1B08",
        x"0B19",
        x"0921",
        x"0931",
        x"2FB3",
        x"2FA2",
        x"2F91",
        x"2F80",
        x"8109",
        x"811A",
        x"812B",
        x"813C",
        x"1B80",
        x"0B91",
        x"0BA2",
        x"0BB3",
        x"2F68",
        x"2F79",
        x"2F8A",
        x"2F9B",
        x"810D",
        x"811E",
        x"812F",
        x"8538",
        x"1B60",
        x"0B71",
        x"0B82",
        x"0B93",
        x"2D23",
        x"E030",
        x"E040",
        x"E050",
        x"940E",
        x"22BC",
        x"2FB5",
        x"2FA4",
        x"2F93",
        x"2F82",
        x"9602",
        x"1DA1",
        x"1DB1",
        x"2DEC",
        x"2DFD",
        x"8F86",
        x"8F97",
        x"A3A0",
        x"A3B1",
        x"3F87",
        x"E0FF",
        x"079F",
        x"05A1",
        x"05B1",
        x"F040",
        x"3F87",
        x"4F9F",
        x"05A1",
        x"05B1",
        x"F008",
        x"C0BD",
        x"E012",
        x"C001",
        x"E011",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"0D84",
        x"1D95",
        x"1DA6",
        x"1DB7",
        x"2DEC",
        x"2DFD",
        x"A386",
        x"A397",
        x"A7A0",
        x"A7B1",
        x"818D",
        x"819E",
        x"81AF",
        x"85B8",
        x"0D84",
        x"1D95",
        x"1DA6",
        x"1DB7",
        x"8129",
        x"813A",
        x"814B",
        x"815C",
        x"0F82",
        x"1F93",
        x"1FA4",
        x"1FB5",
        x"2DEC",
        x"2DFD",
        x"A782",
        x"A793",
        x"A7A4",
        x"A7B5",
        x"EF8F",
        x"EF9F",
        x"EFAF",
        x"EFBF",
        x"8786",
        x"8797",
        x"8BA0",
        x"8BB1",
        x"8214",
        x"3013",
        x"F009",
        x"C05E",
        x"8215",
        x"2DAE",
        x"2DBF",
        x"96D0",
        x"918D",
        x"919C",
        x"97D1",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"0F28",
        x"1F39",
        x"1D41",
        x"1D51",
        x"8B22",
        x"8B33",
        x"8B44",
        x"8B55",
        x"E001",
        x"2D6E",
        x"2D7F",
        x"8181",
        x"940E",
        x"183C",
        x"2B89",
        x"F009",
        x"C042",
        x"2DAC",
        x"2DBD",
        x"96D2",
        x"91ED",
        x"91FC",
        x"97D3",
        x"2FAE",
        x"2FBF",
        x"50A2",
        x"4FBE",
        x"918D",
        x"919C",
        x"3585",
        x"4A9A",
        x"F599",
        x"8180",
        x"8191",
        x"81A2",
        x"81B3",
        x"3582",
        x"4592",
        x"46A1",
        x"44B1",
        x"F551",
        x"2FAE",
        x"2FBF",
        x"51AC",
        x"4FBE",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"3782",
        x"4792",
        x"44A1",
        x"46B1",
        x"F4E1",
        x"2FAE",
        x"2FBF",
        x"51A4",
        x"4FBE",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"2DAC",
        x"2DBD",
        x"961A",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"971D",
        x"51E8",
        x"4FFE",
        x"8180",
        x"8191",
        x"81A2",
        x"81B3",
        x"2DEC",
        x"2DFD",
        x"8786",
        x"8797",
        x"8BA0",
        x"8BB1",
        x"2DAC",
        x"2DBD",
        x"931C",
        x"2DEC",
        x"2DFD",
        x"A616",
        x"A617",
        x"AA10",
        x"AA11",
        x"9656",
        x"921D",
        x"921D",
        x"921D",
        x"921C",
        x"9759",
        x"9180",
        x"009F",
        x"9190",
        x"00A0",
        x"9601",
        x"9390",
        x"00A0",
        x"9380",
        x"009F",
        x"9617",
        x"939C",
        x"938E",
        x"9716",
        x"C006",
        x"E08B",
        x"E090",
        x"C01A",
        x"E08C",
        x"E090",
        x"C017",
        x"E080",
        x"E090",
        x"C014",
        x"E083",
        x"E090",
        x"C011",
        x"E081",
        x"E090",
        x"C00E",
        x"2DEE",
        x"2DFF",
        x"A584",
        x"A595",
        x"A5A6",
        x"A5B7",
        x"2DEC",
        x"2DFD",
        x"A386",
        x"A397",
        x"A7A0",
        x"A7B1",
        x"E013",
        x"CF46",
        x"9628",
        x"E1E1",
        x"940C",
        x"2326",
        x"2388",
        x"F4A1",
        x"91E0",
        x"00A1",
        x"91F0",
        x"00A2",
        x"9730",
        x"F009",
        x"8210",
        x"1561",
        x"0571",
        x"F019",
        x"2FE6",
        x"2FF7",
        x"8210",
        x"9370",
        x"00A2",
        x"9360",
        x"00A1",
        x"E080",
        x"E090",
        x"9508",
        x"E08B",
        x"E090",
        x"9508",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"972E",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2EE8",
        x"2EF9",
        x"877E",
        x"876D",
        x"2EB4",
        x"2FA8",
        x"2FB9",
        x"921D",
        x"921C",
        x"714E",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"0A0F",
        x"9700",
        x"F009",
        x"C121",
        x"2DBB",
        x"71BF",
        x"2EDB",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07FD",
        x"2D2B",
        x"712C",
        x"F409",
        x"C091",
        x"9700",
        x"F099",
        x"3084",
        x"0591",
        x"F009",
        x"C107",
        x"EA88",
        x"E093",
        x"940E",
        x"0973",
        x"9700",
        x"F009",
        x"C100",
        x"2DED",
        x"60E8",
        x"2EDE",
        x"9100",
        x"03BA",
        x"9110",
        x"03BB",
        x"C064",
        x"FCB2",
        x"C0F4",
        x"9100",
        x"03BA",
        x"9110",
        x"03BB",
        x"1501",
        x"0511",
        x"F409",
        x"C0F2",
        x"2FA0",
        x"2FB1",
        x"961B",
        x"918C",
        x"971B",
        x"7181",
        x"F009",
        x"C0EA",
        x"FEB3",
        x"C050",
        x"9654",
        x"908D",
        x"909C",
        x"9755",
        x"2CA1",
        x"2CB1",
        x"2DA8",
        x"2DB9",
        x"2799",
        x"2788",
        x"2FE0",
        x"2FF1",
        x"8C82",
        x"8C93",
        x"2CA1",
        x"2CB1",
        x"2A88",
        x"2A99",
        x"2AAA",
        x"2ABB",
        x"8A15",
        x"8A14",
        x"8E13",
        x"8E12",
        x"8E14",
        x"8E15",
        x"8E16",
        x"8E17",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"E021",
        x"2FE8",
        x"2FF9",
        x"8324",
        x"A446",
        x"A457",
        x"A860",
        x"A871",
        x"1481",
        x"0491",
        x"04A1",
        x"04B1",
        x"F0B1",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"940E",
        x"0551",
        x"9700",
        x"F009",
        x"C0AE",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"E081",
        x"1A88",
        x"0891",
        x"08A1",
        x"08B1",
        x"8682",
        x"8693",
        x"86A4",
        x"86B5",
        x"2D77",
        x"2D66",
        x"2D55",
        x"2D44",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"014C",
        x"9700",
        x"F009",
        x"C094",
        x"FED3",
        x"C02B",
        x"2FA0",
        x"2FB1",
        x"961B",
        x"921C",
        x"940E",
        x"1831",
        x"2FE0",
        x"2FF1",
        x"8766",
        x"8777",
        x"8B80",
        x"8B91",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"E081",
        x"8384",
        x"2DFD",
        x"62F0",
        x"2EDF",
        x"C015",
        x"9700",
        x"F009",
        x"C079",
        x"9100",
        x"03BA",
        x"9110",
        x"03BB",
        x"1501",
        x"0511",
        x"F409",
        x"C073",
        x"2FA0",
        x"2FB1",
        x"961B",
        x"918C",
        x"FD84",
        x"C06D",
        x"FEB1",
        x"C002",
        x"FD80",
        x"C06B",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"A546",
        x"A557",
        x"A960",
        x"A971",
        x"2DAE",
        x"2DBF",
        x"965A",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"975D",
        x"9180",
        x"03BA",
        x"9190",
        x"03BB",
        x"965F",
        x"939C",
        x"938E",
        x"975E",
        x"9614",
        x"92DC",
        x"2FA0",
        x"2FB1",
        x"9654",
        x"918D",
        x"919C",
        x"9755",
        x"E0A0",
        x"E0B0",
        x"2EA8",
        x"2EB9",
        x"2499",
        x"2488",
        x"2FA0",
        x"2FB1",
        x"965A",
        x"914D",
        x"915C",
        x"975B",
        x"E060",
        x"E070",
        x"2948",
        x"2959",
        x"296A",
        x"297B",
        x"2DAE",
        x"2DBF",
        x"961E",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9751",
        x"2FA0",
        x"2FB1",
        x"965C",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"975F",
        x"2DAE",
        x"2DBF",
        x"961A",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"971D",
        x"9616",
        x"921D",
        x"921D",
        x"921D",
        x"921C",
        x"9719",
        x"EF8F",
        x"9615",
        x"938C",
        x"9715",
        x"9656",
        x"921D",
        x"921D",
        x"921D",
        x"921C",
        x"9759",
        x"9611",
        x"93FC",
        x"93EE",
        x"8186",
        x"8197",
        x"9613",
        x"939C",
        x"938E",
        x"9712",
        x"E020",
        x"C007",
        x"E028",
        x"C005",
        x"2F28",
        x"C004",
        x"E024",
        x"C001",
        x"E027",
        x"E090",
        x"2F82",
        x"962E",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"9508",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"839C",
        x"838B",
        x"2EA6",
        x"2EB7",
        x"2EC4",
        x"2ED5",
        x"833A",
        x"8329",
        x"2FA2",
        x"2FB3",
        x"921D",
        x"921C",
        x"2FE8",
        x"2FF9",
        x"8162",
        x"8173",
        x"8180",
        x"8191",
        x"940E",
        x"01FA",
        x"9700",
        x"F009",
        x"C18D",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"FD87",
        x"C182",
        x"FF80",
        x"C182",
        x"961A",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"81EB",
        x"81FC",
        x"8146",
        x"8157",
        x"8560",
        x"8571",
        x"1B84",
        x"0B95",
        x"0BA6",
        x"0BB7",
        x"2D4C",
        x"2D5D",
        x"E060",
        x"E070",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F410",
        x"2EC8",
        x"2ED9",
        x"802B",
        x"803C",
        x"E2F0",
        x"0E2F",
        x"1C31",
        x"14C1",
        x"04D1",
        x"F409",
        x"C15A",
        x"81AB",
        x"81BC",
        x"9616",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9719",
        x"2FB7",
        x"2FA6",
        x"2F95",
        x"2F84",
        x"7091",
        x"27AA",
        x"27BB",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F009",
        x"C105",
        x"81EB",
        x"81FC",
        x"8180",
        x"8191",
        x"8135",
        x"2FA8",
        x"2FB9",
        x"9612",
        x"912C",
        x"1732",
        x"F160",
        x"2B45",
        x"2B46",
        x"2B47",
        x"F429",
        x"8566",
        x"8577",
        x"8980",
        x"8991",
        x"C008",
        x"81EB",
        x"81FC",
        x"8942",
        x"8953",
        x"8964",
        x"8975",
        x"940E",
        x"0282",
        x"3062",
        x"0571",
        x"0581",
        x"0591",
        x"F138",
        x"3F6F",
        x"EFBF",
        x"077B",
        x"078B",
        x"079B",
        x"F431",
        x"81EB",
        x"81FC",
        x"8184",
        x"6880",
        x"8384",
        x"C0CD",
        x"81AB",
        x"81BC",
        x"9652",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"9755",
        x"9615",
        x"921C",
        x"81EB",
        x"81FC",
        x"8080",
        x"8091",
        x"8942",
        x"8953",
        x"8964",
        x"8975",
        x"2D88",
        x"2D99",
        x"940E",
        x"05C4",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F449",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"6880",
        x"9614",
        x"938C",
        x"C0F7",
        x"81EB",
        x"81FC",
        x"8125",
        x"2E46",
        x"2E57",
        x"2E68",
        x"2E79",
        x"0E42",
        x"1C51",
        x"1C61",
        x"1C71",
        x"2CEC",
        x"2CFD",
        x"2CEF",
        x"24FF",
        x"94E6",
        x"14E1",
        x"04F1",
        x"F409",
        x"C054",
        x"2DA8",
        x"2DB9",
        x"9612",
        x"918C",
        x"E030",
        x"2D4E",
        x"2D5F",
        x"0F42",
        x"1F53",
        x"E090",
        x"1784",
        x"0795",
        x"F420",
        x"2EE8",
        x"2EF9",
        x"1AE2",
        x"0AF3",
        x"2D0E",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D6A",
        x"2D7B",
        x"2DE8",
        x"2DF9",
        x"8181",
        x"940E",
        x"183C",
        x"81AB",
        x"81BC",
        x"9614",
        x"912C",
        x"9714",
        x"2B89",
        x"F021",
        x"6820",
        x"9614",
        x"932C",
        x"C06D",
        x"FF26",
        x"C01E",
        x"81EB",
        x"81FC",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1984",
        x"0995",
        x"09A6",
        x"09B7",
        x"2D4E",
        x"2D5F",
        x"E060",
        x"E070",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F458",
        x"2F98",
        x"2788",
        x"0F99",
        x"E040",
        x"E052",
        x"2D62",
        x"2D73",
        x"0D8A",
        x"1D9B",
        x"940E",
        x"00BC",
        x"81AB",
        x"81BC",
        x"9615",
        x"918C",
        x"9715",
        x"0D8E",
        x"9615",
        x"938C",
        x"2CFE",
        x"24EE",
        x"0CFF",
        x"C071",
        x"81EB",
        x"81FC",
        x"8184",
        x"FF86",
        x"C01A",
        x"8926",
        x"8937",
        x"8D40",
        x"8D51",
        x"E001",
        x"2D62",
        x"2D73",
        x"2DA8",
        x"2DB9",
        x"9611",
        x"918C",
        x"940E",
        x"1846",
        x"81EB",
        x"81FC",
        x"8124",
        x"2B89",
        x"F019",
        x"6820",
        x"8324",
        x"C027",
        x"7B2F",
        x"81AB",
        x"81BC",
        x"9614",
        x"932C",
        x"81EB",
        x"81FC",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1584",
        x"0595",
        x"05A6",
        x"05B7",
        x"F0C9",
        x"9001",
        x"81F0",
        x"2DE0",
        x"E001",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D62",
        x"2D73",
        x"8181",
        x"940E",
        x"183C",
        x"2B89",
        x"F051",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"6880",
        x"9614",
        x"938C",
        x"E081",
        x"C04F",
        x"81EB",
        x"81FC",
        x"8A46",
        x"8A57",
        x"8E60",
        x"8E71",
        x"8185",
        x"5F8F",
        x"8385",
        x"81AB",
        x"81BC",
        x"9616",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9719",
        x"2F84",
        x"2F95",
        x"7091",
        x"E0E0",
        x"E0F2",
        x"1BE8",
        x"0BF9",
        x"2CEC",
        x"2CFD",
        x"15EC",
        x"05FD",
        x"F410",
        x"2EEE",
        x"2EFF",
        x"7051",
        x"2766",
        x"2777",
        x"5E40",
        x"4F5F",
        x"816B",
        x"817C",
        x"0F64",
        x"1F75",
        x"2D4E",
        x"2D5F",
        x"2D8A",
        x"2D9B",
        x"940E",
        x"00BC",
        x"0CAE",
        x"1CBF",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"0D8E",
        x"1D9F",
        x"1DA1",
        x"1DB1",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"81A9",
        x"81BA",
        x"918D",
        x"919C",
        x"9711",
        x"0D8E",
        x"1D9F",
        x"938D",
        x"939C",
        x"18CE",
        x"08DF",
        x"CEA2",
        x"E080",
        x"C003",
        x"E082",
        x"C001",
        x"E087",
        x"E090",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"903F",
        x"902F",
        x"9508",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"839C",
        x"838B",
        x"2EA6",
        x"2EB7",
        x"2EC4",
        x"2ED5",
        x"833A",
        x"8329",
        x"2FA2",
        x"2FB3",
        x"921D",
        x"921C",
        x"2FE8",
        x"2FF9",
        x"8162",
        x"8173",
        x"8180",
        x"8191",
        x"940E",
        x"01FA",
        x"9700",
        x"F009",
        x"C1DD",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"FD87",
        x"C1D2",
        x"FF81",
        x"C1D2",
        x"961A",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"0D4C",
        x"1D5D",
        x"1D61",
        x"1D71",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F410",
        x"2CC1",
        x"2CD1",
        x"802B",
        x"803C",
        x"E2B0",
        x"0E2B",
        x"1C31",
        x"14C1",
        x"04D1",
        x"F409",
        x"C04D",
        x"81EB",
        x"81FC",
        x"8146",
        x"8157",
        x"8560",
        x"8571",
        x"2FB7",
        x"2FA6",
        x"2F95",
        x"2F84",
        x"7091",
        x"27AA",
        x"27BB",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F009",
        x"C153",
        x"9001",
        x"81F0",
        x"2DE0",
        x"81AB",
        x"81BC",
        x"9615",
        x"913C",
        x"9715",
        x"8122",
        x"1732",
        x"F408",
        x"C06A",
        x"2B45",
        x"2B46",
        x"2B47",
        x"F4D1",
        x"961E",
        x"916D",
        x"917D",
        x"918D",
        x"919C",
        x"9751",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F5B9",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F8E",
        x"2F9F",
        x"940E",
        x"0469",
        x"81EB",
        x"81FC",
        x"8766",
        x"8777",
        x"8B80",
        x"8B91",
        x"C00C",
        x"81AB",
        x"81BC",
        x"9652",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9755",
        x"2F8E",
        x"2F9F",
        x"940E",
        x"0469",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F4B9",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"8542",
        x"8553",
        x"8564",
        x"8575",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C14B",
        x"81EB",
        x"81FC",
        x"8782",
        x"8793",
        x"87A4",
        x"87B5",
        x"C144",
        x"81AB",
        x"81BC",
        x"9614",
        x"912C",
        x"9714",
        x"3061",
        x"0571",
        x"0581",
        x"0591",
        x"F429",
        x"2F82",
        x"6880",
        x"9614",
        x"938C",
        x"C13F",
        x"3F6F",
        x"EFBF",
        x"077B",
        x"078B",
        x"079B",
        x"F429",
        x"2F82",
        x"6880",
        x"81EB",
        x"81FC",
        x"C0D6",
        x"81AB",
        x"81BC",
        x"9652",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"9755",
        x"9615",
        x"921C",
        x"81EB",
        x"81FC",
        x"8184",
        x"FF86",
        x"C01C",
        x"8926",
        x"8937",
        x"8D40",
        x"8D51",
        x"9001",
        x"81F0",
        x"2DE0",
        x"E001",
        x"2D62",
        x"2D73",
        x"8181",
        x"940E",
        x"1846",
        x"81AB",
        x"81BC",
        x"9614",
        x"912C",
        x"9714",
        x"2B89",
        x"F021",
        x"6820",
        x"9614",
        x"932C",
        x"C0B0",
        x"7B2F",
        x"81EB",
        x"81FC",
        x"8324",
        x"81AB",
        x"81BC",
        x"908D",
        x"909C",
        x"9711",
        x"9652",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9755",
        x"2D88",
        x"2D99",
        x"940E",
        x"05C4",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F431",
        x"81EB",
        x"81FC",
        x"8184",
        x"6880",
        x"8384",
        x"C0EF",
        x"81AB",
        x"81BC",
        x"9615",
        x"912C",
        x"2E46",
        x"2E57",
        x"2E68",
        x"2E79",
        x"0E42",
        x"1C51",
        x"1C61",
        x"1C71",
        x"2CEC",
        x"2CFD",
        x"2CEF",
        x"24FF",
        x"94E6",
        x"14E1",
        x"04F1",
        x"F409",
        x"C051",
        x"2DE8",
        x"2DF9",
        x"8182",
        x"E030",
        x"2D4E",
        x"2D5F",
        x"0F42",
        x"1F53",
        x"E090",
        x"1784",
        x"0795",
        x"F420",
        x"2EE8",
        x"2EF9",
        x"1AE2",
        x"0AF3",
        x"2D0E",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D6A",
        x"2D7B",
        x"2DA8",
        x"2DB9",
        x"9611",
        x"918C",
        x"940E",
        x"1846",
        x"81EB",
        x"81FC",
        x"2B89",
        x"F009",
        x"C058",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1984",
        x"0995",
        x"09A6",
        x"09B7",
        x"2D4E",
        x"2D5F",
        x"E060",
        x"E070",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F4A8",
        x"2F98",
        x"2788",
        x"0F99",
        x"2D6A",
        x"2D7B",
        x"0F68",
        x"1F79",
        x"E040",
        x"E052",
        x"2D82",
        x"2D93",
        x"940E",
        x"00BC",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"7B8F",
        x"9614",
        x"938C",
        x"81EB",
        x"81FC",
        x"8185",
        x"0D8E",
        x"8385",
        x"2CFE",
        x"24EE",
        x"0CFF",
        x"C063",
        x"81EB",
        x"81FC",
        x"8986",
        x"8997",
        x"8DA0",
        x"8DB1",
        x"1584",
        x"0595",
        x"05A6",
        x"05B7",
        x"F119",
        x"8146",
        x"8157",
        x"8560",
        x"8571",
        x"8582",
        x"8593",
        x"85A4",
        x"85B5",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F4B0",
        x"E001",
        x"2D57",
        x"2D46",
        x"2D35",
        x"2D24",
        x"2D62",
        x"2D73",
        x"2DA8",
        x"2DB9",
        x"9611",
        x"918C",
        x"940E",
        x"183C",
        x"2B89",
        x"F039",
        x"81EB",
        x"81FC",
        x"8184",
        x"6880",
        x"8384",
        x"E081",
        x"C05E",
        x"81AB",
        x"81BC",
        x"9656",
        x"924D",
        x"925D",
        x"926D",
        x"927C",
        x"9759",
        x"9615",
        x"918C",
        x"9715",
        x"5F8F",
        x"9615",
        x"938C",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"2F28",
        x"2F39",
        x"7031",
        x"E040",
        x"E052",
        x"1B42",
        x"0B53",
        x"2CEC",
        x"2CFD",
        x"154C",
        x"055D",
        x"F410",
        x"2EE4",
        x"2EF5",
        x"7091",
        x"27AA",
        x"27BB",
        x"9680",
        x"2D4E",
        x"2D5F",
        x"2D6A",
        x"2D7B",
        x"81AB",
        x"81BC",
        x"0F8A",
        x"1F9B",
        x"940E",
        x"00BC",
        x"81EB",
        x"81FC",
        x"8184",
        x"6480",
        x"8384",
        x"0CAE",
        x"1CBF",
        x"81EB",
        x"81FC",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"0D8E",
        x"1D9F",
        x"1DA1",
        x"1DB1",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"81A9",
        x"81BA",
        x"918D",
        x"919C",
        x"9711",
        x"0D8E",
        x"1D9F",
        x"938D",
        x"939C",
        x"18CE",
        x"08DF",
        x"CE54",
        x"81AB",
        x"81BC",
        x"9614",
        x"918C",
        x"9714",
        x"6280",
        x"9614",
        x"938C",
        x"E080",
        x"C003",
        x"E082",
        x"C001",
        x"E087",
        x"E090",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"903F",
        x"902F",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"816A",
        x"817B",
        x"8188",
        x"8199",
        x"940E",
        x"01FA",
        x"9700",
        x"F009",
        x"C051",
        x"818C",
        x"FF85",
        x"C04A",
        x"FF86",
        x"C013",
        x"892E",
        x"893F",
        x"8D48",
        x"8D59",
        x"81E8",
        x"81F9",
        x"E001",
        x"2F6C",
        x"2F7D",
        x"5E60",
        x"4F7F",
        x"8181",
        x"940E",
        x"1846",
        x"2B89",
        x"F5D1",
        x"818C",
        x"7B8F",
        x"838C",
        x"8D4A",
        x"8D5B",
        x"8D6C",
        x"8D7D",
        x"8188",
        x"8199",
        x"940E",
        x"014C",
        x"9700",
        x"F579",
        x"8D0E",
        x"8D1F",
        x"2FE0",
        x"2FF1",
        x"8583",
        x"6280",
        x"8783",
        x"858A",
        x"859B",
        x"85AC",
        x"85BD",
        x"8F84",
        x"8F95",
        x"8FA6",
        x"8FB7",
        x"858E",
        x"859F",
        x"89A8",
        x"89B9",
        x"8F93",
        x"8F82",
        x"8BB5",
        x"8BA4",
        x"940E",
        x"1831",
        x"2FE0",
        x"2FF1",
        x"8B66",
        x"8B77",
        x"8F80",
        x"8F91",
        x"818C",
        x"7D8F",
        x"838C",
        x"81E8",
        x"81F9",
        x"E081",
        x"8384",
        x"8188",
        x"8199",
        x"940E",
        x"0214",
        x"C004",
        x"E080",
        x"C001",
        x"E081",
        x"E090",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"1183",
        x"9700",
        x"F411",
        x"8219",
        x"8218",
        x"91DF",
        x"91CF",
        x"9508",
        x"2388",
        x"F429",
        x"9210",
        x"009E",
        x"E080",
        x"E090",
        x"9508",
        x"E08B",
        x"E090",
        x"9508",
        x"E0AE",
        x"E0B0",
        x"E0E5",
        x"E1F2",
        x"940C",
        x"2317",
        x"879E",
        x"878D",
        x"E040",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"0A0F",
        x"9700",
        x"F009",
        x"C045",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07FD",
        x"9700",
        x"F589",
        x"91A0",
        x"03BA",
        x"91B0",
        x"03BB",
        x"9710",
        x"F449",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"8A16",
        x"8A17",
        x"8E10",
        x"8E11",
        x"C027",
        x"961B",
        x"912C",
        x"971B",
        x"FF24",
        x"C020",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"9654",
        x"914D",
        x"915C",
        x"9755",
        x"E060",
        x"E070",
        x"2F64",
        x"2F75",
        x"2755",
        x"2744",
        x"965A",
        x"910D",
        x"911C",
        x"975B",
        x"E020",
        x"E030",
        x"2B40",
        x"2B51",
        x"2B62",
        x"2B73",
        x"8B46",
        x"8B57",
        x"8F60",
        x"8F71",
        x"C005",
        x"3084",
        x"0591",
        x"F411",
        x"E085",
        x"E090",
        x"962E",
        x"E0E4",
        x"940C",
        x"2333",
        x"E0A4",
        x"E0B0",
        x"E6E1",
        x"E1F2",
        x"940C",
        x"2309",
        x"2E28",
        x"2E39",
        x"2EC4",
        x"2ED5",
        x"2EE6",
        x"2EF7",
        x"2FA8",
        x"2FB9",
        x"9612",
        x"916D",
        x"917C",
        x"9713",
        x"918D",
        x"919C",
        x"940E",
        x"01FA",
        x"9700",
        x"F009",
        x"C1DB",
        x"2DE2",
        x"2DF3",
        x"8124",
        x"FD27",
        x"C1D2",
        x"8582",
        x"8593",
        x"85A4",
        x"85B5",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F430",
        x"FD21",
        x"C004",
        x"2EC8",
        x"2ED9",
        x"2EEA",
        x"2EFB",
        x"2DA2",
        x"2DB3",
        x"9616",
        x"904D",
        x"905D",
        x"906D",
        x"907C",
        x"9719",
        x"2DE2",
        x"2DF3",
        x"8216",
        x"8217",
        x"8610",
        x"8611",
        x"EF8F",
        x"8385",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F429",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"C13D",
        x"8100",
        x"8111",
        x"2FE0",
        x"2FF1",
        x"8082",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"E099",
        x"0C88",
        x"1C99",
        x"1CAA",
        x"1CBB",
        x"959A",
        x"F7D1",
        x"1441",
        x"0451",
        x"0461",
        x"0471",
        x"F409",
        x"C049",
        x"E0F1",
        x"1A4F",
        x"0851",
        x"0861",
        x"0871",
        x"2D9F",
        x"2D8E",
        x"2D7D",
        x"2D6C",
        x"5061",
        x"0971",
        x"0981",
        x"0991",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"940E",
        x"22BC",
        x"8329",
        x"833A",
        x"834B",
        x"835C",
        x"2D97",
        x"2D86",
        x"2D75",
        x"2D64",
        x"2D5B",
        x"2D4A",
        x"2D39",
        x"2D28",
        x"940E",
        x"22BC",
        x"8169",
        x"817A",
        x"818B",
        x"819C",
        x"1762",
        x"0773",
        x"0784",
        x"0795",
        x"F0F8",
        x"2788",
        x"2799",
        x"27AA",
        x"27BB",
        x"1988",
        x"0999",
        x"09AA",
        x"09BB",
        x"2248",
        x"2259",
        x"226A",
        x"227B",
        x"2DA2",
        x"2DB3",
        x"9616",
        x"924D",
        x"925D",
        x"926D",
        x"927C",
        x"9719",
        x"18C4",
        x"08D5",
        x"08E6",
        x"08F7",
        x"9652",
        x"914D",
        x"915D",
        x"916D",
        x"917C",
        x"9755",
        x"C03A",
        x"2DE2",
        x"2DF3",
        x"8546",
        x"8557",
        x"8960",
        x"8971",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F549",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"0469",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"3041",
        x"0551",
        x"0561",
        x"0571",
        x"F449",
        x"2DA2",
        x"2DB3",
        x"9614",
        x"918C",
        x"9714",
        x"6880",
        x"9614",
        x"938C",
        x"C126",
        x"3F4F",
        x"EFBF",
        x"075B",
        x"076B",
        x"077B",
        x"F409",
        x"C0F9",
        x"2DA2",
        x"2DB3",
        x"961E",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9751",
        x"2DE2",
        x"2DF3",
        x"8B42",
        x"8B53",
        x"8B64",
        x"8B75",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F409",
        x"CF5D",
        x"148C",
        x"049D",
        x"04AE",
        x"04BF",
        x"F008",
        x"C057",
        x"2DA2",
        x"2DB3",
        x"9614",
        x"912C",
        x"9714",
        x"918D",
        x"919C",
        x"FF21",
        x"C00C",
        x"940E",
        x"0469",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F439",
        x"C03E",
        x"940E",
        x"0282",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"3F4F",
        x"EFBF",
        x"075B",
        x"076B",
        x"077B",
        x"F409",
        x"C0BD",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F408",
        x"C05E",
        x"2DA2",
        x"2DB3",
        x"91ED",
        x"91FC",
        x"8D86",
        x"8D97",
        x"A1A0",
        x"A1B1",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F008",
        x"C050",
        x"2DA2",
        x"2DB3",
        x"9652",
        x"934D",
        x"935D",
        x"936D",
        x"937C",
        x"9755",
        x"9616",
        x"918D",
        x"919D",
        x"900D",
        x"91BC",
        x"2DA0",
        x"0D88",
        x"1D99",
        x"1DAA",
        x"1DBB",
        x"2DE2",
        x"2DF3",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"18C8",
        x"08D9",
        x"08EA",
        x"08FB",
        x"CFA7",
        x"2CFB",
        x"2CEA",
        x"2CD9",
        x"2CC8",
        x"2DE2",
        x"2DF3",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"0D8C",
        x"1D9D",
        x"1DAE",
        x"1DBF",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"2C8C",
        x"2C9D",
        x"2CAE",
        x"2CBF",
        x"E089",
        x"94B6",
        x"94A7",
        x"9497",
        x"9487",
        x"958A",
        x"F7D1",
        x"8285",
        x"E0F1",
        x"22DF",
        x"24EE",
        x"24FF",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F409",
        x"CEDC",
        x"2DA2",
        x"2DB3",
        x"918D",
        x"919C",
        x"940E",
        x"05C4",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F431",
        x"2DE2",
        x"2DF3",
        x"8184",
        x"6880",
        x"8384",
        x"C079",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"0CC8",
        x"1CD9",
        x"1CEA",
        x"1CFB",
        x"9483",
        x"2DA2",
        x"2DB3",
        x"9615",
        x"928C",
        x"2DE2",
        x"2DF3",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"7091",
        x"27AA",
        x"27BB",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F409",
        x"C047",
        x"8926",
        x"8937",
        x"8D40",
        x"8D51",
        x"16C2",
        x"06D3",
        x"06E4",
        x"06F5",
        x"F1F1",
        x"8184",
        x"2D62",
        x"2D73",
        x"5E60",
        x"4F7F",
        x"2EA6",
        x"2EB7",
        x"FF86",
        x"C016",
        x"9001",
        x"81F0",
        x"2DE0",
        x"E001",
        x"8181",
        x"940E",
        x"1846",
        x"2DA2",
        x"2DB3",
        x"9614",
        x"912C",
        x"9714",
        x"2B89",
        x"F021",
        x"6820",
        x"9614",
        x"932C",
        x"C019",
        x"7B2F",
        x"2DE2",
        x"2DF3",
        x"8324",
        x"2DA2",
        x"2DB3",
        x"91ED",
        x"91FC",
        x"E001",
        x"2D5F",
        x"2D4E",
        x"2D3D",
        x"2D2C",
        x"2D6A",
        x"2D7B",
        x"8181",
        x"940E",
        x"183C",
        x"2B89",
        x"F039",
        x"2DE2",
        x"2DF3",
        x"8184",
        x"6880",
        x"8384",
        x"E081",
        x"C022",
        x"2DA2",
        x"2DB3",
        x"9656",
        x"92CD",
        x"92DD",
        x"92ED",
        x"92FC",
        x"9759",
        x"2DE2",
        x"2DF3",
        x"8186",
        x"8197",
        x"85A0",
        x"85B1",
        x"8542",
        x"8553",
        x"8564",
        x"8575",
        x"1748",
        x"0759",
        x"076A",
        x"077B",
        x"F450",
        x"8782",
        x"8793",
        x"87A4",
        x"87B5",
        x"8184",
        x"6280",
        x"8384",
        x"C002",
        x"E082",
        x"C001",
        x"E080",
        x"E090",
        x"9624",
        x"E1E2",
        x"940C",
        x"2325",
        x"E0AE",
        x"E0B0",
        x"E5E9",
        x"E1F4",
        x"940C",
        x"2317",
        x"2F08",
        x"2F19",
        x"877E",
        x"876D",
        x"E040",
        x"2F68",
        x"2F79",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"0A0F",
        x"9700",
        x"F009",
        x"C049",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2FA0",
        x"2FB1",
        x"9655",
        x"939C",
        x"938E",
        x"9754",
        x"856D",
        x"857E",
        x"2F80",
        x"2F91",
        x"940E",
        x"07FD",
        x"9700",
        x"F5A9",
        x"2FA0",
        x"2FB1",
        x"9652",
        x"91ED",
        x"91FC",
        x"9753",
        x"9730",
        x"F0E1",
        x"8583",
        x"FD84",
        x"C003",
        x"E085",
        x"E090",
        x"C02A",
        x"8984",
        x"8995",
        x"E0A0",
        x"E0B0",
        x"2FA8",
        x"2FB9",
        x"2799",
        x"2788",
        x"8D42",
        x"8D53",
        x"E060",
        x"E070",
        x"2B84",
        x"2B95",
        x"2BA6",
        x"2BB7",
        x"2FE0",
        x"2FF1",
        x"8386",
        x"8397",
        x"87A0",
        x"87B1",
        x"2FA0",
        x"2FB1",
        x"91ED",
        x"91FC",
        x"9711",
        x"8186",
        x"8197",
        x"9613",
        x"939C",
        x"938E",
        x"9712",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"060C",
        x"3084",
        x"0591",
        x"F299",
        x"962E",
        x"E0E4",
        x"940C",
        x"2333",
        x"E0AC",
        x"E0B0",
        x"EBEB",
        x"E1F4",
        x"940C",
        x"2313",
        x"2F08",
        x"2F19",
        x"2EC6",
        x"2ED7",
        x"2FE8",
        x"2FF9",
        x"8162",
        x"8173",
        x"8180",
        x"8191",
        x"940E",
        x"01FA",
        x"2EE8",
        x"2EF9",
        x"2B89",
        x"F5C9",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2FE0",
        x"2FF1",
        x"8B95",
        x"8B84",
        x"14C1",
        x"04D1",
        x"F439",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"060C",
        x"C026",
        x"2F80",
        x"2F91",
        x"940E",
        x"09D0",
        x"3084",
        x"0591",
        x"F439",
        x"2FE0",
        x"2FF1",
        x"8616",
        x"8617",
        x"8A10",
        x"8A11",
        x"C002",
        x"9700",
        x"F4B1",
        x"2D6C",
        x"2D7D",
        x"2F80",
        x"2F91",
        x"940E",
        x"00CB",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"06EB",
        x"3084",
        x"0591",
        x"F439",
        x"2FE0",
        x"2FF1",
        x"8616",
        x"8617",
        x"8A10",
        x"8A11",
        x"C002",
        x"2EE8",
        x"2EF9",
        x"2D8E",
        x"2D9F",
        x"962C",
        x"E0E8",
        x"940C",
        x"232F",
        x"E0AE",
        x"E0B0",
        x"E1E0",
        x"E1F5",
        x"940C",
        x"2315",
        x"879E",
        x"878D",
        x"2EE6",
        x"2EF7",
        x"E040",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"0A0F",
        x"2F08",
        x"2F19",
        x"2B89",
        x"F501",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07FD",
        x"2F08",
        x"2F19",
        x"2B89",
        x"F479",
        x"9180",
        x"03BA",
        x"9190",
        x"03BB",
        x"2B89",
        x"F039",
        x"2D6E",
        x"2D7F",
        x"EA88",
        x"E093",
        x"940E",
        x"00CB",
        x"C002",
        x"E006",
        x"E010",
        x"2F80",
        x"2F91",
        x"962E",
        x"E0E6",
        x"940C",
        x"2331",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"97A4",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"A39C",
        x"A38B",
        x"E041",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"9683",
        x"940E",
        x"0A0F",
        x"9700",
        x"F009",
        x"C083",
        x"2F8C",
        x"2F9D",
        x"9647",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"A16B",
        x"A17C",
        x"EA88",
        x"E093",
        x"940E",
        x"07FD",
        x"9700",
        x"F009",
        x"C073",
        x"91E0",
        x"03BC",
        x"91F0",
        x"03BD",
        x"8583",
        x"FD85",
        x"C06A",
        x"91E0",
        x"03BA",
        x"91F0",
        x"03BB",
        x"9730",
        x"F409",
        x"C060",
        x"8523",
        x"FF20",
        x"C002",
        x"E027",
        x"C05C",
        x"88C4",
        x"88D5",
        x"2CE1",
        x"2CF1",
        x"2CEC",
        x"2CFD",
        x"24DD",
        x"24CC",
        x"8D82",
        x"8D93",
        x"E0A0",
        x"E0B0",
        x"2AC8",
        x"2AD9",
        x"2AEA",
        x"2AFB",
        x"FD24",
        x"C007",
        x"EA88",
        x"E093",
        x"940E",
        x"06CC",
        x"9700",
        x"F141",
        x"C047",
        x"E082",
        x"16C8",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F1D0",
        x"E146",
        x"E050",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"00BC",
        x"82CF",
        x"86D8",
        x"86E9",
        x"86FA",
        x"E062",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"060C",
        x"9700",
        x"F559",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"09D0",
        x"9700",
        x"F211",
        x"3084",
        x"0591",
        x"F299",
        x"C020",
        x"14C1",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F439",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"0214",
        x"C014",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"0551",
        x"9700",
        x"F441",
        x"CFEC",
        x"E022",
        x"C001",
        x"E026",
        x"E090",
        x"C003",
        x"E086",
        x"E090",
        x"2F28",
        x"2F82",
        x"96A4",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"9508",
        x"E1A6",
        x"E0B0",
        x"EFE9",
        x"E1F5",
        x"940C",
        x"2309",
        x"879E",
        x"878D",
        x"E041",
        x"EA68",
        x"E073",
        x"2F8C",
        x"2F9D",
        x"960D",
        x"940E",
        x"0A0F",
        x"9700",
        x"F5A1",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"9390",
        x"03BD",
        x"9380",
        x"03BC",
        x"856D",
        x"857E",
        x"EA88",
        x"E093",
        x"940E",
        x"07FD",
        x"9700",
        x"F069",
        x"3084",
        x"0591",
        x"F511",
        x"91E0",
        x"03BC",
        x"91F0",
        x"03BD",
        x"8583",
        x"FF85",
        x"C01D",
        x"E086",
        x"E090",
        x"C018",
        x"E088",
        x"E090",
        x"C015",
        x"91E0",
        x"03BA",
        x"91F0",
        x"03BB",
        x"E120",
        x"8723",
        x"8A46",
        x"8A57",
        x"8E60",
        x"8E71",
        x"8ED3",
        x"8EC2",
        x"8A95",
        x"8A84",
        x"E021",
        x"2FA8",
        x"2FB9",
        x"9614",
        x"932C",
        x"940E",
        x"0214",
        x"2F28",
        x"C0FD",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"0469",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"2B67",
        x"2B68",
        x"2B69",
        x"F041",
        x"E031",
        x"16C3",
        x"04D1",
        x"04E1",
        x"04F1",
        x"F421",
        x"E022",
        x"C009",
        x"E027",
        x"C007",
        x"EFBF",
        x"16CB",
        x"06DB",
        x"06EB",
        x"06FB",
        x"F419",
        x"E021",
        x"E090",
        x"C0D8",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"940E",
        x"014C",
        x"9700",
        x"F669",
        x"9100",
        x"03A8",
        x"9110",
        x"03A9",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2F80",
        x"2F91",
        x"940E",
        x"05C4",
        x"8B6B",
        x"877F",
        x"2F38",
        x"8B9C",
        x"2FA0",
        x"2FB1",
        x"96D2",
        x"910D",
        x"911C",
        x"97D3",
        x"2E20",
        x"2E31",
        x"EFBE",
        x"1A3B",
        x"2FE0",
        x"2FF1",
        x"15E2",
        x"05F3",
        x"F011",
        x"9211",
        x"CFFB",
        x"2F80",
        x"2F91",
        x"960B",
        x"2FE0",
        x"2FF1",
        x"E240",
        x"17E8",
        x"07F9",
        x"F011",
        x"9341",
        x"CFFB",
        x"E22E",
        x"2FE0",
        x"2FF1",
        x"8320",
        x"E180",
        x"8783",
        x"8B2E",
        x"8B3D",
        x"940E",
        x"1831",
        x"2E46",
        x"2E57",
        x"2E68",
        x"2E79",
        x"2FA0",
        x"2FB1",
        x"9656",
        x"936D",
        x"937D",
        x"938D",
        x"939C",
        x"9759",
        x"965B",
        x"92DC",
        x"92CE",
        x"975A",
        x"2C9F",
        x"2C8E",
        x"24AA",
        x"24BB",
        x"9655",
        x"929C",
        x"928E",
        x"9754",
        x"E240",
        x"E050",
        x"2F60",
        x"2F71",
        x"2F80",
        x"2F91",
        x"9680",
        x"940E",
        x"00BC",
        x"892E",
        x"2FE0",
        x"2FF1",
        x"A321",
        x"9180",
        x"03AE",
        x"9190",
        x"03AF",
        x"91A0",
        x"03B0",
        x"91B0",
        x"03B1",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"8140",
        x"893D",
        x"3043",
        x"F469",
        x"A146",
        x"A157",
        x"A560",
        x"A571",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F421",
        x"E080",
        x"E090",
        x"E0A0",
        x"E0B0",
        x"2FE0",
        x"2FF1",
        x"AF93",
        x"AF82",
        x"ABB5",
        x"ABA4",
        x"894B",
        x"855F",
        x"2F63",
        x"897C",
        x"E021",
        x"91E0",
        x"03A8",
        x"91F0",
        x"03A9",
        x"8192",
        x"2F84",
        x"893B",
        x"1B83",
        x"1789",
        x"F548",
        x"2FB7",
        x"2FA6",
        x"2F95",
        x"2F84",
        x"9601",
        x"1DA1",
        x"1DB1",
        x"878F",
        x"8B98",
        x"8BA9",
        x"8BBA",
        x"A746",
        x"A757",
        x"AB60",
        x"AB71",
        x"8324",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F8E",
        x"2F9F",
        x"8B2E",
        x"940E",
        x"014C",
        x"892E",
        x"9700",
        x"F009",
        x"CF23",
        x"2FE0",
        x"2FF1",
        x"15E2",
        x"05F3",
        x"F011",
        x"9211",
        x"CFFB",
        x"854F",
        x"8958",
        x"8969",
        x"897A",
        x"CFCD",
        x"EA88",
        x"E093",
        x"940E",
        x"0973",
        x"2F08",
        x"2F19",
        x"9180",
        x"03A8",
        x"9190",
        x"03A9",
        x"1501",
        x"0511",
        x"F409",
        x"CEF4",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"940E",
        x"0551",
        x"2F20",
        x"2F91",
        x"2F82",
        x"9666",
        x"E1E2",
        x"940C",
        x"2325",
        x"E4AF",
        x"E0B0",
        x"E4E3",
        x"E1F7",
        x"940C",
        x"2315",
        x"9660",
        x"AF9F",
        x"AF8E",
        x"9760",
        x"2F06",
        x"2F17",
        x"2F8C",
        x"2F9D",
        x"5B8E",
        x"4F9F",
        x"A79C",
        x"A78B",
        x"E041",
        x"2F6C",
        x"2F7D",
        x"5E69",
        x"4F7F",
        x"960C",
        x"940E",
        x"0A0F",
        x"9700",
        x"F009",
        x"C0D0",
        x"898F",
        x"8D98",
        x"839A",
        x"8389",
        x"9660",
        x"AD6E",
        x"AD7F",
        x"9760",
        x"2F8C",
        x"2F9D",
        x"9647",
        x"940E",
        x"07FD",
        x"9700",
        x"F009",
        x"C0C0",
        x"A5EB",
        x"A5FC",
        x"8583",
        x"FD85",
        x"C0AA",
        x"A589",
        x"A59A",
        x"9700",
        x"F409",
        x"C0A2",
        x"2F68",
        x"2F79",
        x"5F65",
        x"4F7F",
        x"E145",
        x"E050",
        x"2F8C",
        x"2F9D",
        x"968D",
        x"940E",
        x"00BC",
        x"E146",
        x"E050",
        x"2F6C",
        x"2F7D",
        x"5E69",
        x"4F7F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"00BC",
        x"2F60",
        x"2F71",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"07FD",
        x"9700",
        x"F409",
        x"C080",
        x"3084",
        x"0591",
        x"F009",
        x"C092",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"0973",
        x"9700",
        x"F009",
        x"C08A",
        x"88EB",
        x"88FC",
        x"E143",
        x"E050",
        x"2F6C",
        x"2F7D",
        x"5D61",
        x"4F7F",
        x"2D8E",
        x"2D9F",
        x"960D",
        x"940E",
        x"00BC",
        x"A58D",
        x"6280",
        x"2DAE",
        x"2DBF",
        x"961B",
        x"938C",
        x"971B",
        x"89EF",
        x"8DF8",
        x"E081",
        x"8384",
        x"961B",
        x"918C",
        x"971B",
        x"FF84",
        x"C05F",
        x"8109",
        x"811A",
        x"965A",
        x"914D",
        x"915C",
        x"975B",
        x"9654",
        x"912D",
        x"913C",
        x"9755",
        x"2B42",
        x"2B53",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"05C4",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"1541",
        x"0551",
        x"0561",
        x"0571",
        x"F409",
        x"C04F",
        x"2F80",
        x"2F91",
        x"940E",
        x"014C",
        x"81E9",
        x"81FA",
        x"A922",
        x"A933",
        x"9700",
        x"F009",
        x"C046",
        x"2FA2",
        x"2FB3",
        x"9691",
        x"918C",
        x"328E",
        x"F591",
        x"8140",
        x"818F",
        x"8598",
        x"85A9",
        x"85BA",
        x"3043",
        x"F449",
        x"A146",
        x"A157",
        x"A560",
        x"A571",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F029",
        x"2F78",
        x"2F69",
        x"2F5A",
        x"2F4B",
        x"C004",
        x"E070",
        x"E060",
        x"E050",
        x"E040",
        x"2F87",
        x"2F96",
        x"2FA2",
        x"2FB3",
        x"96DB",
        x"939C",
        x"938E",
        x"97DA",
        x"2F85",
        x"2F94",
        x"96D5",
        x"939C",
        x"938E",
        x"97D4",
        x"E081",
        x"8384",
        x"C008",
        x"E028",
        x"C001",
        x"E024",
        x"E090",
        x"C012",
        x"E086",
        x"E090",
        x"C00E",
        x"2F8C",
        x"2F9D",
        x"9647",
        x"940E",
        x"06CC",
        x"9700",
        x"F439",
        x"898F",
        x"8D98",
        x"940E",
        x"0214",
        x"C002",
        x"E082",
        x"E090",
        x"2F28",
        x"2F82",
        x"5BC1",
        x"4FDF",
        x"E0E6",
        x"940C",
        x"2331",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"9508",
        x"940E",
        x"18B6",
        x"9508",
        x"940E",
        x"18AE",
        x"9508",
        x"2F86",
        x"2F97",
        x"2F75",
        x"2F64",
        x"2F53",
        x"2F42",
        x"940E",
        x"1957",
        x"E090",
        x"9508",
        x"2F86",
        x"2F97",
        x"2F75",
        x"2F64",
        x"2F53",
        x"2F42",
        x"940E",
        x"19F8",
        x"E090",
        x"9508",
        x"E080",
        x"E090",
        x"9508",
        x"B381",
        x"6B80",
        x"BB81",
        x"988E",
        x"9A6C",
        x"B18D",
        x"7F8C",
        x"B98D",
        x"9A6E",
        x"9A94",
        x"9A97",
        x"9508",
        x"B98F",
        x"9B77",
        x"CFFE",
        x"B18F",
        x"9508",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD4",
        x"2F15",
        x"2F06",
        x"2EF7",
        x"FF87",
        x"C00A",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E787",
        x"940E",
        x"1864",
        x"3082",
        x"F558",
        x"77CF",
        x"9A94",
        x"EF8F",
        x"940E",
        x"185F",
        x"9894",
        x"EF8F",
        x"940E",
        x"185F",
        x"2F8C",
        x"940E",
        x"185F",
        x"2D8F",
        x"940E",
        x"185F",
        x"2F80",
        x"940E",
        x"185F",
        x"2F81",
        x"940E",
        x"185F",
        x"2F8D",
        x"940E",
        x"185F",
        x"34C0",
        x"F021",
        x"34C8",
        x"F421",
        x"E887",
        x"C003",
        x"E985",
        x"C001",
        x"E081",
        x"940E",
        x"185F",
        x"E0CA",
        x"EF8F",
        x"940E",
        x"185F",
        x"FF87",
        x"C002",
        x"50C1",
        x"F7C9",
        x"B7CD",
        x"B7DE",
        x"E0E5",
        x"940C",
        x"2332",
        x"9A94",
        x"EF8F",
        x"940E",
        x"185F",
        x"9508",
        x"9180",
        x"03BE",
        x"2388",
        x"F011",
        x"E080",
        x"9508",
        x"E082",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"EBEC",
        x"E1F8",
        x"940C",
        x"2314",
        x"98C6",
        x"940E",
        x"1853",
        x"E01B",
        x"EF8F",
        x"940E",
        x"185F",
        x"5011",
        x"F7D9",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E480",
        x"940E",
        x"1864",
        x"3081",
        x"F009",
        x"C082",
        x"EA4A",
        x"E051",
        x"E060",
        x"E070",
        x"E488",
        x"940E",
        x"1864",
        x"3081",
        x"F569",
        x"2F0C",
        x"2F1D",
        x"5F0F",
        x"4F1F",
        x"2EE0",
        x"2EF1",
        x"E024",
        x"2ED2",
        x"0ED0",
        x"EF8F",
        x"940E",
        x"185F",
        x"2DEE",
        x"2DFF",
        x"9381",
        x"2EEE",
        x"2EFF",
        x"16DE",
        x"F7B1",
        x"818B",
        x"3081",
        x"F009",
        x"C062",
        x"818C",
        x"3A8A",
        x"F009",
        x"C05E",
        x"EE90",
        x"2EE9",
        x"E29E",
        x"2EF9",
        x"E040",
        x"E050",
        x"E060",
        x"E470",
        x"EE89",
        x"940E",
        x"1864",
        x"2388",
        x"F129",
        x"E0F1",
        x"1AEF",
        x"08F1",
        x"F799",
        x"C04C",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"EE89",
        x"940E",
        x"1864",
        x"3082",
        x"F018",
        x"E011",
        x"E401",
        x"C002",
        x"E012",
        x"EE09",
        x"EA88",
        x"2EE8",
        x"E681",
        x"2EF8",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"2F80",
        x"940E",
        x"1864",
        x"2388",
        x"F141",
        x"E0F1",
        x"1AEF",
        x"08F1",
        x"F799",
        x"C02C",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E78A",
        x"940E",
        x"1864",
        x"2388",
        x"F519",
        x"EF8F",
        x"940E",
        x"185F",
        x"2FE0",
        x"2FF1",
        x"9381",
        x"2F0E",
        x"2F1F",
        x"16DE",
        x"F7B1",
        x"8189",
        x"FD86",
        x"C002",
        x"E014",
        x"C001",
        x"E01C",
        x"9310",
        x"03BE",
        x"940E",
        x"18A9",
        x"9AC6",
        x"E081",
        x"2311",
        x"F069",
        x"E080",
        x"C00B",
        x"E040",
        x"E052",
        x"E060",
        x"E070",
        x"E580",
        x"940E",
        x"1864",
        x"2388",
        x"F369",
        x"E010",
        x"CFEB",
        x"9624",
        x"E0E7",
        x"940C",
        x"2330",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"98C6",
        x"9180",
        x"03BE",
        x"FD83",
        x"C007",
        x"E089",
        x"0F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"958A",
        x"F7D1",
        x"E581",
        x"940E",
        x"1864",
        x"2388",
        x"F019",
        x"E0C1",
        x"E0D0",
        x"C020",
        x"E3C0",
        x"E7D5",
        x"EF8F",
        x"940E",
        x"185F",
        x"3F8F",
        x"F419",
        x"9721",
        x"F7C9",
        x"CFF3",
        x"3F8E",
        x"F789",
        x"2FC0",
        x"2FD1",
        x"2F0C",
        x"2F1D",
        x"5F1E",
        x"EF8F",
        x"940E",
        x"185F",
        x"9389",
        x"17C0",
        x"07D1",
        x"F7C9",
        x"EF8F",
        x"940E",
        x"185F",
        x"EF8F",
        x"940E",
        x"185F",
        x"E0C0",
        x"E0D0",
        x"940E",
        x"18A9",
        x"9AC6",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"92EF",
        x"92FF",
        x"931F",
        x"93CF",
        x"93DF",
        x"2EF8",
        x"2EE9",
        x"2F12",
        x"98C6",
        x"9180",
        x"03BE",
        x"FD83",
        x"C007",
        x"E089",
        x"0F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"958A",
        x"F7D1",
        x"E581",
        x"940E",
        x"1864",
        x"2388",
        x"F019",
        x"E0C1",
        x"E0D0",
        x"C036",
        x"E3C0",
        x"E7D5",
        x"EF8F",
        x"940E",
        x"185F",
        x"3F8F",
        x"F419",
        x"9721",
        x"F7C9",
        x"CFF3",
        x"3F8E",
        x"F789",
        x"2311",
        x"F431",
        x"2DCF",
        x"2DDE",
        x"2EEC",
        x"2EFD",
        x"94F3",
        x"C008",
        x"E0C0",
        x"E0D1",
        x"EF8F",
        x"940E",
        x"185F",
        x"9721",
        x"F7D9",
        x"CFF2",
        x"EF8F",
        x"940E",
        x"185F",
        x"9389",
        x"15CE",
        x"05DF",
        x"F7C9",
        x"2311",
        x"F049",
        x"EF8F",
        x"940E",
        x"185F",
        x"EF8F",
        x"940E",
        x"185F",
        x"E0C0",
        x"E0D0",
        x"C008",
        x"E0C0",
        x"E0D1",
        x"EF8F",
        x"940E",
        x"185F",
        x"9721",
        x"F7D9",
        x"CFEF",
        x"940E",
        x"18A9",
        x"9AC6",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"911F",
        x"90FF",
        x"90EF",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"EFEE",
        x"E1F9",
        x"940C",
        x"2315",
        x"2F08",
        x"2F19",
        x"98C6",
        x"9180",
        x"03BE",
        x"FD83",
        x"C007",
        x"E089",
        x"0F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"958A",
        x"F7D1",
        x"E588",
        x"940E",
        x"1864",
        x"2388",
        x"F019",
        x"E081",
        x"E090",
        x"C03D",
        x"EF8F",
        x"940E",
        x"185F",
        x"EF8E",
        x"940E",
        x"185F",
        x"2EE0",
        x"2EF1",
        x"2D0E",
        x"2D1F",
        x"5F1E",
        x"2DEE",
        x"2DFF",
        x"9181",
        x"2EEE",
        x"2EFF",
        x"940E",
        x"185F",
        x"16E0",
        x"06F1",
        x"F7B1",
        x"E080",
        x"940E",
        x"185F",
        x"E080",
        x"940E",
        x"185F",
        x"EF8F",
        x"940E",
        x"185F",
        x"718F",
        x"3085",
        x"F6E1",
        x"EE08",
        x"EF1D",
        x"EF8F",
        x"940E",
        x"185F",
        x"3F8F",
        x"F049",
        x"1501",
        x"0511",
        x"F019",
        x"5001",
        x"0911",
        x"CFF5",
        x"E081",
        x"E090",
        x"C006",
        x"E081",
        x"E090",
        x"1501",
        x"0511",
        x"F009",
        x"E080",
        x"8389",
        x"839A",
        x"940E",
        x"18A9",
        x"819A",
        x"8189",
        x"9AC6",
        x"9622",
        x"E0E6",
        x"940C",
        x"2331",
        x"93CF",
        x"93DF",
        x"9AC3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"0000",
        x"B389",
        x"9380",
        x"00A3",
        x"9AC0",
        x"9180",
        x"00A3",
        x"2F98",
        x"7190",
        x"FD84",
        x"C002",
        x"9380",
        x"00A4",
        x"9180",
        x"00A4",
        x"7087",
        x"3081",
        x"F409",
        x"C176",
        x"F038",
        x"3082",
        x"F409",
        x"C143",
        x"3083",
        x"F409",
        x"C153",
        x"C1CC",
        x"2399",
        x"F009",
        x"C1C9",
        x"98C3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"0000",
        x"B389",
        x"9380",
        x"00A5",
        x"9AC0",
        x"9180",
        x"00A5",
        x"2F98",
        x"7998",
        x"3190",
        x"F451",
        x"2F28",
        x"9522",
        x"9526",
        x"7027",
        x"E030",
        x"9330",
        x"0064",
        x"9320",
        x"0063",
        x"798F",
        x"2F98",
        x"7F90",
        x"3290",
        x"F459",
        x"2F28",
        x"9526",
        x"9526",
        x"7023",
        x"E030",
        x"9330",
        x"0064",
        x"9320",
        x"0063",
        x"7F83",
        x"C006",
        x"2388",
        x"F409",
        x"C15A",
        x"3081",
        x"F409",
        x"C171",
        x"3082",
        x"F409",
        x"C171",
        x"3084",
        x"F409",
        x"C171",
        x"3085",
        x"F409",
        x"C171",
        x"3088",
        x"F409",
        x"C171",
        x"3180",
        x"F409",
        x"C171",
        x"3181",
        x"F409",
        x"C171",
        x"3182",
        x"F409",
        x"C171",
        x"3183",
        x"F409",
        x"C171",
        x"3187",
        x"F409",
        x"C171",
        x"3184",
        x"F409",
        x"C171",
        x"3185",
        x"F409",
        x"C171",
        x"3186",
        x"F409",
        x"C171",
        x"3280",
        x"F481",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"02A8",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"E081",
        x"9380",
        x"03FF",
        x"E082",
        x"9380",
        x"00A4",
        x"C041",
        x"3281",
        x"F429",
        x"9210",
        x"03FF",
        x"9210",
        x"03FA",
        x"C03A",
        x"3282",
        x"F451",
        x"9180",
        x"03BF",
        x"E090",
        x"9390",
        x"046F",
        x"9380",
        x"046E",
        x"E9C5",
        x"E1DE",
        x"C122",
        x"3283",
        x"F451",
        x"9180",
        x"03BF",
        x"E090",
        x"9390",
        x"046F",
        x"9380",
        x"046E",
        x"EEC0",
        x"E1DE",
        x"C116",
        x"338F",
        x"F409",
        x"C140",
        x"3480",
        x"F501",
        x"9180",
        x"02A8",
        x"7083",
        x"9380",
        x"03F9",
        x"9180",
        x"02A9",
        x"9190",
        x"02AA",
        x"91A0",
        x"02AB",
        x"91B0",
        x"02AC",
        x"9380",
        x"03FB",
        x"9390",
        x"03FC",
        x"93A0",
        x"03FD",
        x"93B0",
        x"03FE",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"E0C0",
        x"E0D0",
        x"C0F1",
        x"3481",
        x"F489",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"03BF",
        x"7083",
        x"E090",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"5480",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8585",
        x"C0C5",
        x"E0C0",
        x"E0D0",
        x"3482",
        x"F409",
        x"C0C8",
        x"3483",
        x"F409",
        x"C0C8",
        x"3484",
        x"F409",
        x"C0C8",
        x"3485",
        x"F409",
        x"C0C8",
        x"3486",
        x"F409",
        x"C0C8",
        x"3487",
        x"F409",
        x"C0C8",
        x"3880",
        x"F449",
        x"E080",
        x"940E",
        x"1836",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"03BE",
        x"C04B",
        x"3A80",
        x"F429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"B182",
        x"C044",
        x"3A81",
        x"F421",
        x"9180",
        x"03BF",
        x"B982",
        x"C00C",
        x"3A82",
        x"F429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"B181",
        x"C037",
        x"3A83",
        x"F441",
        x"9180",
        x"03BF",
        x"B983",
        x"9160",
        x"03BF",
        x"EF8E",
        x"E090",
        x"C01F",
        x"3E80",
        x"F429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E28C",
        x"C026",
        x"3E81",
        x"F431",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"02A6",
        x"C01E",
        x"3F80",
        x"F431",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"02A7",
        x"C016",
        x"3F81",
        x"F469",
        x"9160",
        x"03BF",
        x"9360",
        x"02A7",
        x"EF8F",
        x"E090",
        x"940E",
        x"23CB",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"C007",
        x"3F8D",
        x"F451",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"00A4",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"C06F",
        x"3F8E",
        x"F009",
        x"C06C",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0060",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9180",
        x"0060",
        x"9580",
        x"9380",
        x"0060",
        x"C05D",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"91E0",
        x"03FF",
        x"E0F0",
        x"55E8",
        x"4FFD",
        x"8180",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9180",
        x"03FF",
        x"5F8F",
        x"9380",
        x"03FF",
        x"C07A",
        x"2399",
        x"F009",
        x"C077",
        x"98C3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"0000",
        x"B389",
        x"9380",
        x"00A5",
        x"9AC0",
        x"9180",
        x"03FF",
        x"2FE8",
        x"E0F0",
        x"55E8",
        x"4FFD",
        x"9190",
        x"00A5",
        x"8390",
        x"5F8F",
        x"9380",
        x"03FF",
        x"E081",
        x"9380",
        x"03FA",
        x"C05E",
        x"2399",
        x"F009",
        x"C05B",
        x"98C3",
        x"BA1A",
        x"98C0",
        x"0000",
        x"0000",
        x"B389",
        x"9380",
        x"00A5",
        x"9AC0",
        x"9180",
        x"00A5",
        x"9380",
        x"03BF",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"03BF",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"C044",
        x"E0CD",
        x"E1DD",
        x"C011",
        x"E9C9",
        x"E2D1",
        x"C00E",
        x"E4C6",
        x"E2D0",
        x"C00B",
        x"E9C5",
        x"E2D0",
        x"C008",
        x"E5CF",
        x"E2D1",
        x"C005",
        x"EFC9",
        x"E2D0",
        x"C002",
        x"E6CA",
        x"E2D1",
        x"9720",
        x"F171",
        x"2FEC",
        x"2FFD",
        x"9509",
        x"C02A",
        x"E2C8",
        x"E1DD",
        x"CFF7",
        x"E9CC",
        x"E1DD",
        x"CFF4",
        x"EAC9",
        x"E1DD",
        x"CFF1",
        x"EBC6",
        x"E1DD",
        x"CFEE",
        x"ECC3",
        x"E1DD",
        x"CFEB",
        x"E1C4",
        x"E1DF",
        x"CFE8",
        x"EDC7",
        x"E1DD",
        x"CFE5",
        x"EFC8",
        x"E1DF",
        x"CFE2",
        x"EFC6",
        x"E1DD",
        x"CFDF",
        x"E0C2",
        x"E1DE",
        x"CFDC",
        x"E2C9",
        x"E1DF",
        x"CFD9",
        x"E0CE",
        x"E1DE",
        x"CFD6",
        x"E3C6",
        x"E1DF",
        x"CFD3",
        x"EDC4",
        x"E2D1",
        x"CFD0",
        x"91DF",
        x"91CF",
        x"9508",
        x"2F48",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"2B89",
        x"F439",
        x"EA68",
        x"E072",
        x"E780",
        x"E094",
        x"940E",
        x"0C2C",
        x"C03D",
        x"9210",
        x"0064",
        x"9210",
        x"0063",
        x"9180",
        x"0690",
        x"9190",
        x"0691",
        x"2B89",
        x"F419",
        x"E081",
        x"E090",
        x"C011",
        x"9180",
        x"08B0",
        x"9190",
        x"08B1",
        x"2B89",
        x"F419",
        x"E082",
        x"E090",
        x"C008",
        x"9180",
        x"0AD0",
        x"9190",
        x"0AD1",
        x"2B89",
        x"F431",
        x"E083",
        x"E090",
        x"9390",
        x"0064",
        x"9380",
        x"0063",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"1618",
        x"0619",
        x"F494",
        x"E260",
        x"E072",
        x"940E",
        x"22AB",
        x"EA68",
        x"E072",
        x"5980",
        x"4F9B",
        x"940E",
        x"0C2C",
        x"9700",
        x"F441",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"6280",
        x"C002",
        x"E182",
        x"E090",
        x"6480",
        x"9508",
        x"9210",
        x"03F8",
        x"EA86",
        x"E090",
        x"9390",
        x"0D35",
        x"9380",
        x"0D34",
        x"E348",
        x"E050",
        x"EF6F",
        x"E070",
        x"EC80",
        x"E093",
        x"940E",
        x"23A1",
        x"E080",
        x"940E",
        x"11F5",
        x"E062",
        x"E07D",
        x"E080",
        x"940E",
        x"0C13",
        x"9210",
        x"0471",
        x"9210",
        x"0470",
        x"9210",
        x"0691",
        x"9210",
        x"0690",
        x"9210",
        x"08B1",
        x"9210",
        x"08B0",
        x"9210",
        x"0AD1",
        x"9210",
        x"0AD0",
        x"9508",
        x"EAE8",
        x"E0F2",
        x"9001",
        x"2000",
        x"F7E9",
        x"9731",
        x"5AE8",
        x"40F2",
        x"EAA8",
        x"E0B2",
        x"EF6F",
        x"EF7F",
        x"EF2F",
        x"EF3F",
        x"E080",
        x"E090",
        x"178E",
        x"079F",
        x"F139",
        x"3F2F",
        x"EF4F",
        x"0734",
        x"F489",
        x"914D",
        x"334F",
        x"F039",
        x"324A",
        x"F029",
        x"354C",
        x"F031",
        x"324F",
        x"F431",
        x"C003",
        x"2F28",
        x"2F39",
        x"C002",
        x"2F68",
        x"2F79",
        x"9601",
        x"CFE8",
        x"3F6F",
        x"EF8F",
        x"0778",
        x"F0D1",
        x"2FE6",
        x"2FF7",
        x"55E8",
        x"4FFD",
        x"8210",
        x"5567",
        x"4F7D",
        x"E140",
        x"E050",
        x"EF81",
        x"E09C",
        x"940E",
        x"23B2",
        x"9508",
        x"3F2F",
        x"4F3F",
        x"F759",
        x"E140",
        x"E050",
        x"E768",
        x"E070",
        x"EF81",
        x"E09C",
        x"940E",
        x"2380",
        x"9508",
        x"E140",
        x"E050",
        x"EA68",
        x"E072",
        x"EF81",
        x"E09C",
        x"940E",
        x"23B2",
        x"9210",
        x"02A8",
        x"9508",
        x"940E",
        x"1CBC",
        x"EA68",
        x"E072",
        x"E588",
        x"E094",
        x"940E",
        x"1453",
        x"9380",
        x"0CF0",
        x"98C3",
        x"2388",
        x"F031",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0CF0",
        x"6480",
        x"C003",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"E060",
        x"E074",
        x"E588",
        x"E094",
        x"940E",
        x"14B5",
        x"9380",
        x"0CF0",
        x"2388",
        x"F421",
        x"9180",
        x"0409",
        x"2388",
        x"F439",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0CF0",
        x"6480",
        x"C051",
        x"E069",
        x"E074",
        x"EF81",
        x"E09C",
        x"940E",
        x"2234",
        x"2B89",
        x"F319",
        x"E0E9",
        x"E0F4",
        x"9001",
        x"2000",
        x"F7E9",
        x"2F0E",
        x"2F1F",
        x"500A",
        x"4014",
        x"2FC0",
        x"91D0",
        x"0408",
        x"2F8D",
        x"7180",
        x"2EF8",
        x"FFD4",
        x"C005",
        x"E38C",
        x"9380",
        x"02A8",
        x"E081",
        x"C001",
        x"E080",
        x"2E08",
        x"0C00",
        x"0B99",
        x"E069",
        x"E074",
        x"5588",
        x"4F9D",
        x"940E",
        x"23A9",
        x"20FF",
        x"F059",
        x"2FE0",
        x"2E00",
        x"0C00",
        x"0BFF",
        x"55E8",
        x"4FFD",
        x"E38E",
        x"8381",
        x"8212",
        x"E0C2",
        x"0FC0",
        x"2F8C",
        x"0FCC",
        x"0B99",
        x"2FE8",
        x"2FF9",
        x"55E8",
        x"4FFD",
        x"83D1",
        x"2FE8",
        x"2FF9",
        x"55E6",
        x"4FFD",
        x"9140",
        x"0400",
        x"9150",
        x"0401",
        x"9160",
        x"0402",
        x"9170",
        x"0403",
        x"8340",
        x"8351",
        x"8362",
        x"8373",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"B7CD",
        x"B7DE",
        x"E0E5",
        x"940C",
        x"2332",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"11FF",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"15F3",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"1546",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"EAE8",
        x"E0F2",
        x"9001",
        x"2000",
        x"F7E9",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"2F6E",
        x"2F7F",
        x"EA88",
        x"E092",
        x"940E",
        x"173D",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"E081",
        x"940E",
        x"1C46",
        x"9380",
        x"0CF0",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"3084",
        x"0591",
        x"F444",
        x"E166",
        x"E070",
        x"940E",
        x"22AB",
        x"5080",
        x"4F9C",
        x"940E",
        x"0A08",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"9180",
        x"0CF0",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E086",
        x"940E",
        x"1C46",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E182",
        x"940E",
        x"1C46",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E1E4",
        x"E1FE",
        x"940C",
        x"230D",
        x"9100",
        x"0063",
        x"9110",
        x"0064",
        x"2F80",
        x"2F91",
        x"E260",
        x"E072",
        x"940E",
        x"22AB",
        x"5980",
        x"4F9B",
        x"2FE8",
        x"2FF9",
        x"963A",
        x"2FA8",
        x"2FB9",
        x"961A",
        x"913C",
        x"971A",
        x"8121",
        x"8192",
        x"8183",
        x"EAC8",
        x"E0D2",
        x"8338",
        x"8329",
        x"839A",
        x"838B",
        x"E082",
        x"2E68",
        x"E08D",
        x"2E78",
        x"2DE6",
        x"2DF7",
        x"8082",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"2FEA",
        x"2FFB",
        x"8586",
        x"8597",
        x"89A0",
        x"89B1",
        x"2F28",
        x"2F39",
        x"2F4A",
        x"2F5B",
        x"5022",
        x"0931",
        x"0941",
        x"0951",
        x"2D9B",
        x"2D8A",
        x"2D79",
        x"2D68",
        x"940E",
        x"22E5",
        x"2E82",
        x"2E93",
        x"2EA4",
        x"2EB5",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"2DE6",
        x"2DF7",
        x"A582",
        x"A593",
        x"A5A4",
        x"A5B5",
        x"0D88",
        x"1D99",
        x"1DAA",
        x"1DBB",
        x"838C",
        x"839D",
        x"83AE",
        x"83BF",
        x"2F80",
        x"2F91",
        x"E260",
        x"E072",
        x"940E",
        x"22AB",
        x"5980",
        x"4F9B",
        x"2FE8",
        x"2FF9",
        x"9636",
        x"2FA8",
        x"2FB9",
        x"9616",
        x"913C",
        x"8121",
        x"8192",
        x"8183",
        x"8738",
        x"8729",
        x"879A",
        x"878B",
        x"2F80",
        x"2F91",
        x"E166",
        x"E070",
        x"940E",
        x"22AB",
        x"5080",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8580",
        x"738F",
        x"878C",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"B7CD",
        x"B7DE",
        x"E0EE",
        x"940C",
        x"2329",
        x"E0A2",
        x"E0B0",
        x"E9EB",
        x"E1FE",
        x"940C",
        x"2319",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"22AB",
        x"5980",
        x"4F9B",
        x"9120",
        x"046E",
        x"9130",
        x"046F",
        x"2B23",
        x"F431",
        x"E020",
        x"E031",
        x"9330",
        x"046F",
        x"9320",
        x"046E",
        x"9140",
        x"046E",
        x"9150",
        x"046F",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"EA68",
        x"E072",
        x"940E",
        x"0D95",
        x"9120",
        x"0063",
        x"9130",
        x"0064",
        x"1612",
        x"0613",
        x"F484",
        x"9700",
        x"F471",
        x"9140",
        x"046E",
        x"9150",
        x"046F",
        x"8129",
        x"813A",
        x"1742",
        x"0753",
        x"F029",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E680",
        x"C004",
        x"98C3",
        x"EF9F",
        x"BB9A",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"2335",
        x"E0A2",
        x"E0B0",
        x"EEE6",
        x"E1FE",
        x"940C",
        x"2319",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"22AB",
        x"5980",
        x"4F9B",
        x"9120",
        x"046E",
        x"9130",
        x"046F",
        x"2B23",
        x"F431",
        x"E020",
        x"E031",
        x"9330",
        x"046F",
        x"9320",
        x"046E",
        x"98C3",
        x"EF2F",
        x"BB2A",
        x"9140",
        x"046E",
        x"9150",
        x"046F",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"EA68",
        x"E072",
        x"940E",
        x"0F64",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"2335",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"22AB",
        x"98C3",
        x"EF2F",
        x"BB2A",
        x"5980",
        x"4F9B",
        x"940E",
        x"11E8",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"EA88",
        x"E092",
        x"940E",
        x"1546",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"9180",
        x"0063",
        x"9190",
        x"0064",
        x"E260",
        x"E072",
        x"940E",
        x"22AB",
        x"EAE8",
        x"E0F2",
        x"8140",
        x"8151",
        x"8162",
        x"8173",
        x"98C3",
        x"EF2F",
        x"BB2A",
        x"5980",
        x"4F9B",
        x"940E",
        x"125B",
        x"6480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"93CF",
        x"93DF",
        x"9120",
        x"0061",
        x"9130",
        x"0062",
        x"1782",
        x"0793",
        x"F419",
        x"E080",
        x"E090",
        x"C025",
        x"2FC8",
        x"2FD9",
        x"FD37",
        x"C004",
        x"ED80",
        x"E09A",
        x"940E",
        x"11E8",
        x"EF8F",
        x"EF9F",
        x"9390",
        x"0062",
        x"9380",
        x"0061",
        x"FDD7",
        x"CFED",
        x"2F8C",
        x"2F9D",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"2F68",
        x"2F79",
        x"5460",
        x"4F7C",
        x"E043",
        x"ED80",
        x"E09A",
        x"940E",
        x"0C2C",
        x"9700",
        x"F421",
        x"93D0",
        x"0062",
        x"93C0",
        x"0061",
        x"91DF",
        x"91CF",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"940E",
        x"1F51",
        x"9380",
        x"0CF0",
        x"2388",
        x"F019",
        x"2F28",
        x"6420",
        x"C031",
        x"2F80",
        x"2F91",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"5480",
        x"4F9C",
        x"2EE8",
        x"2EF9",
        x"ECC0",
        x"E0D3",
        x"16EC",
        x"06FD",
        x"F051",
        x"E04E",
        x"E050",
        x"2F6C",
        x"2F7D",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"2392",
        x"2B89",
        x"F0B9",
        x"962E",
        x"E083",
        x"3FC8",
        x"07D8",
        x"F771",
        x"E080",
        x"E094",
        x"940E",
        x"0A08",
        x"9120",
        x"0408",
        x"2F80",
        x"2F91",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"5480",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8725",
        x"C001",
        x"E42A",
        x"2F82",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"2331",
        x"E0A2",
        x"E0B0",
        x"EDE3",
        x"E1FF",
        x"940C",
        x"2319",
        x"E66C",
        x"E070",
        x"EA88",
        x"E092",
        x"940E",
        x"2376",
        x"E142",
        x"EA68",
        x"E072",
        x"E780",
        x"E094",
        x"940E",
        x"0C2C",
        x"9380",
        x"0CF0",
        x"2388",
        x"F481",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E348",
        x"E050",
        x"EC60",
        x"E073",
        x"E780",
        x"E094",
        x"940E",
        x"0F64",
        x"E780",
        x"E094",
        x"940E",
        x"11E8",
        x"9622",
        x"E0E2",
        x"940C",
        x"2335",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"91C0",
        x"02A8",
        x"70C3",
        x"E0D0",
        x"2F8C",
        x"2F9D",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"2F08",
        x"2F19",
        x"5400",
        x"4F1C",
        x"E08E",
        x"2FE0",
        x"2FF1",
        x"9211",
        x"958A",
        x"F7E9",
        x"E04D",
        x"E050",
        x"EA69",
        x"E072",
        x"2F80",
        x"2F91",
        x"940E",
        x"23B2",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1F85",
        x"2FC8",
        x"3480",
        x"F040",
        x"E04E",
        x"E050",
        x"EF6F",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"23A1",
        x"940E",
        x"1FCD",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"BBCB",
        x"98C1",
        x"0000",
        x"9AC1",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"9140",
        x"03FB",
        x"9150",
        x"03FC",
        x"9160",
        x"03FD",
        x"9170",
        x"03FE",
        x"2F76",
        x"2F65",
        x"2F54",
        x"2744",
        x"ED80",
        x"E09A",
        x"940E",
        x"125B",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"E4EC",
        x"E2F0",
        x"940C",
        x"2319",
        x"9120",
        x"03F9",
        x"E030",
        x"2F82",
        x"2F93",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"5480",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8585",
        x"3F8F",
        x"F169",
        x"2F82",
        x"2F93",
        x"940E",
        x"1F51",
        x"940E",
        x"2035",
        x"2388",
        x"F4A9",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E040",
        x"E051",
        x"EA68",
        x"E072",
        x"ED80",
        x"E09A",
        x"940E",
        x"0D95",
        x"2F28",
        x"2388",
        x"F439",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"C015",
        x"E429",
        x"9180",
        x"03F9",
        x"E090",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"5480",
        x"4F9C",
        x"EF3F",
        x"2FE8",
        x"2FF9",
        x"8735",
        x"6420",
        x"C001",
        x"E429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"BB2B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"2335",
        x"E0A2",
        x"E0B0",
        x"E9EB",
        x"E2F0",
        x"940C",
        x"2319",
        x"9120",
        x"03F9",
        x"E030",
        x"2F82",
        x"2F93",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"5480",
        x"4F9C",
        x"2FE8",
        x"2FF9",
        x"8585",
        x"3F8F",
        x"F409",
        x"C041",
        x"FF80",
        x"C005",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E48A",
        x"C022",
        x"2F82",
        x"2F93",
        x"940E",
        x"1F51",
        x"940E",
        x"2035",
        x"2388",
        x"F4E1",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E040",
        x"E051",
        x"EA68",
        x"E072",
        x"ED80",
        x"E09A",
        x"940E",
        x"0F64",
        x"2F28",
        x"2388",
        x"F471",
        x"ED80",
        x"E09A",
        x"940E",
        x"1183",
        x"2F28",
        x"2388",
        x"F439",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"C01B",
        x"E429",
        x"9180",
        x"03F9",
        x"E090",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"2FE8",
        x"2FF9",
        x"54E0",
        x"4FFC",
        x"EF9F",
        x"8795",
        x"98C3",
        x"BB9A",
        x"E480",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"C001",
        x"E429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"BB2B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E2",
        x"940C",
        x"2335",
        x"E0A2",
        x"E0B0",
        x"EFEF",
        x"E2F0",
        x"940C",
        x"2313",
        x"E660",
        x"E070",
        x"EA88",
        x"E092",
        x"940E",
        x"2376",
        x"E041",
        x"EA68",
        x"E072",
        x"E780",
        x"E094",
        x"940E",
        x"0C2C",
        x"9380",
        x"0CF0",
        x"2388",
        x"F499",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"E348",
        x"E050",
        x"EC60",
        x"E073",
        x"E780",
        x"E094",
        x"940E",
        x"0D95",
        x"9380",
        x"0CF0",
        x"E780",
        x"E094",
        x"940E",
        x"11E8",
        x"C008",
        x"E348",
        x"E050",
        x"EF6F",
        x"E070",
        x"EC80",
        x"E093",
        x"940E",
        x"23A1",
        x"E000",
        x"E010",
        x"2CE1",
        x"2CF1",
        x"2F80",
        x"2F91",
        x"5480",
        x"4F9C",
        x"2EC8",
        x"2ED9",
        x"2FE8",
        x"2FF9",
        x"8585",
        x"3F8F",
        x"F449",
        x"E04E",
        x"E050",
        x"EF6F",
        x"E070",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"23A1",
        x"C006",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"1F85",
        x"FD86",
        x"CFF1",
        x"EFFF",
        x"1AEF",
        x"0AFF",
        x"5F02",
        x"4F1F",
        x"3308",
        x"0511",
        x"F6F1",
        x"940E",
        x"1FCD",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9622",
        x"E0E8",
        x"940C",
        x"232F",
        x"940E",
        x"1FCD",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"9508",
        x"93CF",
        x"93DF",
        x"91C0",
        x"03BF",
        x"70C3",
        x"E0D0",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1F51",
        x"ED80",
        x"E09A",
        x"940E",
        x"11E8",
        x"EF8F",
        x"EF9F",
        x"9390",
        x"0062",
        x"9380",
        x"0061",
        x"2F8C",
        x"2F9D",
        x"E06E",
        x"E070",
        x"940E",
        x"22AB",
        x"E04E",
        x"E050",
        x"EF6F",
        x"E070",
        x"5480",
        x"4F9C",
        x"940E",
        x"23A1",
        x"940E",
        x"1FCD",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"91DF",
        x"91CF",
        x"9508",
        x"93CF",
        x"93DF",
        x"E020",
        x"E030",
        x"E040",
        x"2FA2",
        x"2FB3",
        x"54A0",
        x"4FBC",
        x"961D",
        x"918C",
        x"971D",
        x"3F8F",
        x"F411",
        x"2FE4",
        x"C014",
        x"E080",
        x"E090",
        x"2FE4",
        x"0FE8",
        x"2FCA",
        x"2FDB",
        x"0FC8",
        x"1FD9",
        x"8158",
        x"2355",
        x"F049",
        x"9601",
        x"308D",
        x"0591",
        x"F029",
        x"E0F0",
        x"55E8",
        x"4FFD",
        x"8350",
        x"CFEE",
        x"2FAE",
        x"E0B0",
        x"55A8",
        x"4FBD",
        x"921C",
        x"E041",
        x"0F4E",
        x"5F22",
        x"4F3F",
        x"3328",
        x"0531",
        x"F6A9",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"91DF",
        x"91CF",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"9180",
        x"046E",
        x"9190",
        x"046F",
        x"2B89",
        x"F449",
        x"9180",
        x"03FA",
        x"2388",
        x"F429",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E488",
        x"C042",
        x"9180",
        x"02A8",
        x"9190",
        x"02A9",
        x"3485",
        x"E522",
        x"0792",
        x"F079",
        x"3485",
        x"4597",
        x"F5D9",
        x"91C0",
        x"02AA",
        x"E0D0",
        x"9180",
        x"02AB",
        x"2EEC",
        x"2EFD",
        x"0EE8",
        x"1CF1",
        x"EA0C",
        x"E012",
        x"C019",
        x"91C0",
        x"02AA",
        x"E0D0",
        x"9180",
        x"02AB",
        x"2EEC",
        x"2EFD",
        x"0EE8",
        x"1CF1",
        x"EA08",
        x"E012",
        x"15CE",
        x"05DF",
        x"F4C8",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"23C3",
        x"2FE0",
        x"2FF1",
        x"9381",
        x"2F0E",
        x"2F1F",
        x"9621",
        x"CFF2",
        x"15CE",
        x"05DF",
        x"F458",
        x"2FE0",
        x"2FF1",
        x"9161",
        x"2F0E",
        x"2F1F",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"23CB",
        x"9621",
        x"CFF2",
        x"98C3",
        x"EF8F",
        x"BB8A",
        x"E38F",
        x"BB8B",
        x"98C1",
        x"0000",
        x"9AC1",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"2331",
        x"93CF",
        x"93DF",
        x"2F28",
        x"2F39",
        x"2FA6",
        x"2FB7",
        x"2FE2",
        x"2FF3",
        x"2FC6",
        x"2FD7",
        x"9189",
        x"2F6C",
        x"2F7D",
        x"2388",
        x"F069",
        x"2FC2",
        x"2FD3",
        x"9199",
        x"2F2C",
        x"2F3D",
        x"329A",
        x"F031",
        x"1798",
        x"F361",
        x"339F",
        x"F351",
        x"E080",
        x"C033",
        x"E040",
        x"E050",
        x"E020",
        x"E030",
        x"919C",
        x"2399",
        x"F111",
        x"8180",
        x"328A",
        x"F469",
        x"2F8E",
        x"2F9F",
        x"9601",
        x"8121",
        x"2322",
        x"F111",
        x"2F2A",
        x"2F3B",
        x"5F2F",
        x"4F3F",
        x"2F48",
        x"2F59",
        x"C00F",
        x"1789",
        x"F011",
        x"338F",
        x"F429",
        x"2F8E",
        x"2F9F",
        x"9601",
        x"9611",
        x"C006",
        x"2FA2",
        x"2FB3",
        x"5F2F",
        x"4F3F",
        x"2F84",
        x"2F95",
        x"2FE8",
        x"2FF9",
        x"CFDB",
        x"9121",
        x"322A",
        x"F3E9",
        x"E081",
        x"E090",
        x"2322",
        x"F021",
        x"E080",
        x"C002",
        x"E081",
        x"E090",
        x"91DF",
        x"91CF",
        x"9508",
        x"E020",
        x"EE31",
        x"E040",
        x"E050",
        x"E060",
        x"EE71",
        x"E080",
        x"E090",
        x"940E",
        x"00B8",
        x"940E",
        x"0087",
        x"9AC7",
        x"9AC6",
        x"B387",
        x"6C80",
        x"BB87",
        x"EF8F",
        x"9380",
        x"02A7",
        x"940E",
        x"1853",
        x"940E",
        x"1C93",
        x"9478",
        x"E180",
        x"BF89",
        x"B608",
        x"FE04",
        x"CFFD",
        x"B788",
        x"6180",
        x"BF88",
        x"940E",
        x"1A56",
        x"CFF7",
        x"2400",
        x"2755",
        x"C004",
        x"0E08",
        x"1F59",
        x"0F88",
        x"1F99",
        x"9700",
        x"F029",
        x"9576",
        x"9567",
        x"F3B8",
        x"0571",
        x"F7B9",
        x"2D80",
        x"2F95",
        x"9508",
        x"E2A1",
        x"2E1A",
        x"1BAA",
        x"1BBB",
        x"2FEA",
        x"2FFB",
        x"C00D",
        x"1FAA",
        x"1FBB",
        x"1FEE",
        x"1FFF",
        x"17A2",
        x"07B3",
        x"07E4",
        x"07F5",
        x"F020",
        x"1BA2",
        x"0BB3",
        x"0BE4",
        x"0BF5",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"941A",
        x"F769",
        x"9560",
        x"9570",
        x"9580",
        x"9590",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"9468",
        x"1300",
        x"94E8",
        x"E0A0",
        x"E0B0",
        x"EEEC",
        x"E2F2",
        x"940C",
        x"2311",
        x"EFEF",
        x"F9E7",
        x"2EA2",
        x"2EB3",
        x"2EC4",
        x"2ED5",
        x"235E",
        x"0F55",
        x"08EE",
        x"2CFE",
        x"2D0E",
        x"2D1F",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"239E",
        x"0F99",
        x"0B66",
        x"2F76",
        x"2F86",
        x"2F97",
        x"940E",
        x"2341",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"232D",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"1BCA",
        x"0BDB",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"9409",
        x"882A",
        x"8839",
        x"8848",
        x"845F",
        x"846E",
        x"847D",
        x"848C",
        x"849B",
        x"84AA",
        x"84B9",
        x"84C8",
        x"80DF",
        x"80EE",
        x"80FD",
        x"810C",
        x"811B",
        x"81AA",
        x"81B9",
        x"0FCE",
        x"1DD1",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2FCA",
        x"2FDB",
        x"9508",
        x"93DF",
        x"93CF",
        x"929F",
        x"E4A0",
        x"2E9A",
        x"2400",
        x"2DA0",
        x"2DB1",
        x"2DC0",
        x"2DD1",
        x"2DE0",
        x"2DF1",
        x"9516",
        x"9507",
        x"94F7",
        x"94E7",
        x"94D7",
        x"94C7",
        x"94B7",
        x"94A7",
        x"F448",
        x"6810",
        x"0FA2",
        x"1FB3",
        x"1FC4",
        x"1FD5",
        x"1FE6",
        x"1FF7",
        x"1E08",
        x"1E19",
        x"0F22",
        x"1F33",
        x"1F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"949A",
        x"F721",
        x"2F2A",
        x"2F3B",
        x"2F4C",
        x"2F5D",
        x"2F6E",
        x"2F7F",
        x"2D80",
        x"2D91",
        x"2411",
        x"909F",
        x"91CF",
        x"91DF",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"95C8",
        x"9631",
        x"920D",
        x"2000",
        x"F7D9",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"5041",
        x"4050",
        x"F050",
        x"95C8",
        x"9631",
        x"920D",
        x"2000",
        x"F7C1",
        x"C001",
        x"921D",
        x"5041",
        x"4050",
        x"F7E0",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"C004",
        x"918D",
        x"9001",
        x"1980",
        x"F421",
        x"5041",
        x"4050",
        x"F7C8",
        x"1B88",
        x"0B99",
        x"9508",
        x"2FA8",
        x"2FB9",
        x"C001",
        x"936D",
        x"5041",
        x"4050",
        x"F7E0",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"9001",
        x"920D",
        x"2000",
        x"F7E1",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"5041",
        x"4050",
        x"F048",
        x"9001",
        x"920D",
        x"2000",
        x"F7C9",
        x"C001",
        x"921D",
        x"5041",
        x"4050",
        x"F7E0",
        x"9508",
        x"99E1",
        x"CFFE",
        x"BB9F",
        x"BB8E",
        x"9AE0",
        x"2799",
        x"B38D",
        x"9508",
        x"2F26",
        x"99E1",
        x"CFFE",
        x"BB9F",
        x"BB8E",
        x"BB2D",
        x"B60F",
        x"94F8",
        x"9AE2",
        x"9AE1",
        x"BE0F",
        x"9601",
        x"9508",
        x"94F8",
        x"CFFF",
        x"FF55",
        x"FFFF",
        x"99FF",
        x"6A21",
        x"5F21",
        x"F921",
        x"9520",
        x"4620",
        x"F820",
        x"D41F",
        x"3621",
        x"291F",
        x"141F",
        x"E01F",
        x"951E",
        x"0E1E",
        x"021E",
        x"F61E",
        x"D71D",
        x"C31D",
        x"B61D",
        x"A91D",
        x"9C1D",
        x"281D",
        x"0D1D",
        x"201D",
        x"2A22",
        x"2C2B",
        x"3D5B",
        x"7C5D",
        x"007F",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF",
        x"FFFF"
    );

begin

    process (cp2)
    begin
        if rising_edge(cp2) then
            if ce = '1' then
                if (we = '1') then
                    RAM(conv_integer(address)) <= din;
                end if;
                dout <= RAM(conv_integer(address));
            end if;
        end if;
    end process;

end RTL;
