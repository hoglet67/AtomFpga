library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity atomfloat is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of atomfloat is

  signal rom_addr : std_logic_vector(11 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(11 downto 0) <= ADDR;
  end process;

  p_rom : process
  begin
    wait until rising_edge(CLK);
    DATA <= (others => '0');
    case rom_addr is
      when x"000" => DATA <= x"AA";
      when x"001" => DATA <= x"55";
      when x"002" => DATA <= x"0E";
      when x"003" => DATA <= x"D1";
      when x"004" => DATA <= x"5E";
      when x"005" => DATA <= x"D1";
      when x"006" => DATA <= x"28";
      when x"007" => DATA <= x"D0";
      when x"008" => DATA <= x"E4";
      when x"009" => DATA <= x"41";
      when x"00A" => DATA <= x"43";
      when x"00B" => DATA <= x"53";
      when x"00C" => DATA <= x"D2";
      when x"00D" => DATA <= x"1E";
      when x"00E" => DATA <= x"41";
      when x"00F" => DATA <= x"53";
      when x"010" => DATA <= x"4E";
      when x"011" => DATA <= x"D2";
      when x"012" => DATA <= x"24";
      when x"013" => DATA <= x"41";
      when x"014" => DATA <= x"54";
      when x"015" => DATA <= x"4E";
      when x"016" => DATA <= x"DC";
      when x"017" => DATA <= x"64";
      when x"018" => DATA <= x"41";
      when x"019" => DATA <= x"42";
      when x"01A" => DATA <= x"53";
      when x"01B" => DATA <= x"D2";
      when x"01C" => DATA <= x"15";
      when x"01D" => DATA <= x"43";
      when x"01E" => DATA <= x"4F";
      when x"01F" => DATA <= x"53";
      when x"020" => DATA <= x"DC";
      when x"021" => DATA <= x"E3";
      when x"022" => DATA <= x"45";
      when x"023" => DATA <= x"58";
      when x"024" => DATA <= x"50";
      when x"025" => DATA <= x"DD";
      when x"026" => DATA <= x"D4";
      when x"027" => DATA <= x"48";
      when x"028" => DATA <= x"54";
      when x"029" => DATA <= x"4E";
      when x"02A" => DATA <= x"DE";
      when x"02B" => DATA <= x"72";
      when x"02C" => DATA <= x"4C";
      when x"02D" => DATA <= x"4F";
      when x"02E" => DATA <= x"47";
      when x"02F" => DATA <= x"DB";
      when x"030" => DATA <= x"B3";
      when x"031" => DATA <= x"50";
      when x"032" => DATA <= x"49";
      when x"033" => DATA <= x"D2";
      when x"034" => DATA <= x"C3";
      when x"035" => DATA <= x"53";
      when x"036" => DATA <= x"49";
      when x"037" => DATA <= x"4E";
      when x"038" => DATA <= x"DC";
      when x"039" => DATA <= x"EE";
      when x"03A" => DATA <= x"53";
      when x"03B" => DATA <= x"51";
      when x"03C" => DATA <= x"52";
      when x"03D" => DATA <= x"DB";
      when x"03E" => DATA <= x"6F";
      when x"03F" => DATA <= x"54";
      when x"040" => DATA <= x"41";
      when x"041" => DATA <= x"4E";
      when x"042" => DATA <= x"DA";
      when x"043" => DATA <= x"C4";
      when x"044" => DATA <= x"44";
      when x"045" => DATA <= x"45";
      when x"046" => DATA <= x"47";
      when x"047" => DATA <= x"D2";
      when x"048" => DATA <= x"73";
      when x"049" => DATA <= x"52";
      when x"04A" => DATA <= x"41";
      when x"04B" => DATA <= x"44";
      when x"04C" => DATA <= x"D2";
      when x"04D" => DATA <= x"65";
      when x"04E" => DATA <= x"53";
      when x"04F" => DATA <= x"47";
      when x"050" => DATA <= x"4E";
      when x"051" => DATA <= x"D2";
      when x"052" => DATA <= x"86";
      when x"053" => DATA <= x"56";
      when x"054" => DATA <= x"41";
      when x"055" => DATA <= x"4C";
      when x"056" => DATA <= x"D2";
      when x"057" => DATA <= x"E0";
      when x"058" => DATA <= x"46";
      when x"059" => DATA <= x"4C";
      when x"05A" => DATA <= x"54";
      when x"05B" => DATA <= x"D2";
      when x"05C" => DATA <= x"9A";
      when x"05D" => DATA <= x"46";
      when x"05E" => DATA <= x"47";
      when x"05F" => DATA <= x"45";
      when x"060" => DATA <= x"54";
      when x"061" => DATA <= x"D2";
      when x"062" => DATA <= x"CC";
      when x"063" => DATA <= x"D2";
      when x"064" => DATA <= x"96";
      when x"065" => DATA <= x"25";
      when x"066" => DATA <= x"D3";
      when x"067" => DATA <= x"0B";
      when x"068" => DATA <= x"46";
      when x"069" => DATA <= x"49";
      when x"06A" => DATA <= x"46";
      when x"06B" => DATA <= x"D3";
      when x"06C" => DATA <= x"A8";
      when x"06D" => DATA <= x"46";
      when x"06E" => DATA <= x"55";
      when x"06F" => DATA <= x"4E";
      when x"070" => DATA <= x"54";
      when x"071" => DATA <= x"49";
      when x"072" => DATA <= x"4C";
      when x"073" => DATA <= x"D3";
      when x"074" => DATA <= x"AE";
      when x"075" => DATA <= x"43";
      when x"076" => DATA <= x"4F";
      when x"077" => DATA <= x"4C";
      when x"078" => DATA <= x"4F";
      when x"079" => DATA <= x"55";
      when x"07A" => DATA <= x"52";
      when x"07B" => DATA <= x"DF";
      when x"07C" => DATA <= x"02";
      when x"07D" => DATA <= x"46";
      when x"07E" => DATA <= x"44";
      when x"07F" => DATA <= x"49";
      when x"080" => DATA <= x"4D";
      when x"081" => DATA <= x"D3";
      when x"082" => DATA <= x"D3";
      when x"083" => DATA <= x"53";
      when x"084" => DATA <= x"54";
      when x"085" => DATA <= x"52";
      when x"086" => DATA <= x"D3";
      when x"087" => DATA <= x"1F";
      when x"088" => DATA <= x"46";
      when x"089" => DATA <= x"50";
      when x"08A" => DATA <= x"52";
      when x"08B" => DATA <= x"49";
      when x"08C" => DATA <= x"4E";
      when x"08D" => DATA <= x"54";
      when x"08E" => DATA <= x"D3";
      when x"08F" => DATA <= x"31";
      when x"090" => DATA <= x"46";
      when x"091" => DATA <= x"49";
      when x"092" => DATA <= x"4E";
      when x"093" => DATA <= x"50";
      when x"094" => DATA <= x"55";
      when x"095" => DATA <= x"54";
      when x"096" => DATA <= x"D3";
      when x"097" => DATA <= x"6A";
      when x"098" => DATA <= x"46";
      when x"099" => DATA <= x"50";
      when x"09A" => DATA <= x"55";
      when x"09B" => DATA <= x"54";
      when x"09C" => DATA <= x"D3";
      when x"09D" => DATA <= x"B4";
      when x"09E" => DATA <= x"D4";
      when x"09F" => DATA <= x"AF";
      when x"0A0" => DATA <= x"2B";
      when x"0A1" => DATA <= x"D1";
      when x"0A2" => DATA <= x"77";
      when x"0A3" => DATA <= x"2D";
      when x"0A4" => DATA <= x"D1";
      when x"0A5" => DATA <= x"83";
      when x"0A6" => DATA <= x"FE";
      when x"0A7" => DATA <= x"2A";
      when x"0A8" => DATA <= x"D1";
      when x"0A9" => DATA <= x"8F";
      when x"0AA" => DATA <= x"2F";
      when x"0AB" => DATA <= x"D1";
      when x"0AC" => DATA <= x"9B";
      when x"0AD" => DATA <= x"FE";
      when x"0AE" => DATA <= x"5E";
      when x"0AF" => DATA <= x"D1";
      when x"0B0" => DATA <= x"A7";
      when x"0B1" => DATA <= x"FE";
      when x"0B2" => DATA <= x"2B";
      when x"0B3" => DATA <= x"D1";
      when x"0B4" => DATA <= x"CB";
      when x"0B5" => DATA <= x"2D";
      when x"0B6" => DATA <= x"D1";
      when x"0B7" => DATA <= x"BC";
      when x"0B8" => DATA <= x"D1";
      when x"0B9" => DATA <= x"CB";
      when x"0BA" => DATA <= x"29";
      when x"0BB" => DATA <= x"C2";
      when x"0BC" => DATA <= x"78";
      when x"0BD" => DATA <= x"FF";
      when x"0BE" => DATA <= x"3B";
      when x"0BF" => DATA <= x"C5";
      when x"0C0" => DATA <= x"4A";
      when x"0C1" => DATA <= x"0D";
      when x"0C2" => DATA <= x"C5";
      when x"0C3" => DATA <= x"4A";
      when x"0C4" => DATA <= x"2C";
      when x"0C5" => DATA <= x"D3";
      when x"0C6" => DATA <= x"31";
      when x"0C7" => DATA <= x"D3";
      when x"0C8" => DATA <= x"39";
      when x"0C9" => DATA <= x"2C";
      when x"0CA" => DATA <= x"D3";
      when x"0CB" => DATA <= x"6A";
      when x"0CC" => DATA <= x"C5";
      when x"0CD" => DATA <= x"58";
      when x"0CE" => DATA <= x"3D";
      when x"0CF" => DATA <= x"D9";
      when x"0D0" => DATA <= x"F6";
      when x"0D1" => DATA <= x"3C";
      when x"0D2" => DATA <= x"3E";
      when x"0D3" => DATA <= x"D9";
      when x"0D4" => DATA <= x"FE";
      when x"0D5" => DATA <= x"3C";
      when x"0D6" => DATA <= x"3D";
      when x"0D7" => DATA <= x"D9";
      when x"0D8" => DATA <= x"FA";
      when x"0D9" => DATA <= x"3C";
      when x"0DA" => DATA <= x"DA";
      when x"0DB" => DATA <= x"02";
      when x"0DC" => DATA <= x"3E";
      when x"0DD" => DATA <= x"3D";
      when x"0DE" => DATA <= x"DA";
      when x"0DF" => DATA <= x"06";
      when x"0E0" => DATA <= x"3E";
      when x"0E1" => DATA <= x"DA";
      when x"0E2" => DATA <= x"0A";
      when x"0E3" => DATA <= x"FF";
      when x"0E4" => DATA <= x"20";
      when x"0E5" => DATA <= x"FC";
      when x"0E6" => DATA <= x"D0";
      when x"0E7" => DATA <= x"A2";
      when x"0E8" => DATA <= x"B4";
      when x"0E9" => DATA <= x"D0";
      when x"0EA" => DATA <= x"20";
      when x"0EB" => DATA <= x"18";
      when x"0EC" => DATA <= x"66";
      when x"0ED" => DATA <= x"73";
      when x"0EE" => DATA <= x"A2";
      when x"0EF" => DATA <= x"AC";
      when x"0F0" => DATA <= x"D0";
      when x"0F1" => DATA <= x"19";
      when x"0F2" => DATA <= x"20";
      when x"0F3" => DATA <= x"5D";
      when x"0F4" => DATA <= x"D8";
      when x"0F5" => DATA <= x"20";
      when x"0F6" => DATA <= x"06";
      when x"0F7" => DATA <= x"D1";
      when x"0F8" => DATA <= x"A2";
      when x"0F9" => DATA <= x"A1";
      when x"0FA" => DATA <= x"D0";
      when x"0FB" => DATA <= x"0F";
      when x"0FC" => DATA <= x"20";
      when x"0FD" => DATA <= x"F5";
      when x"0FE" => DATA <= x"D0";
      when x"0FF" => DATA <= x"A2";
      when x"100" => DATA <= x"9A";
      when x"101" => DATA <= x"D0";
      when x"102" => DATA <= x"08";
      when x"103" => DATA <= x"20";
      when x"104" => DATA <= x"5D";
      when x"105" => DATA <= x"D8";
      when x"106" => DATA <= x"20";
      when x"107" => DATA <= x"EB";
      when x"108" => DATA <= x"D0";
      when x"109" => DATA <= x"A2";
      when x"10A" => DATA <= x"A8";
      when x"10B" => DATA <= x"18";
      when x"10C" => DATA <= x"90";
      when x"10D" => DATA <= x"05";
      when x"10E" => DATA <= x"A2";
      when x"10F" => DATA <= x"5F";
      when x"110" => DATA <= x"84";
      when x"111" => DATA <= x"03";
      when x"112" => DATA <= x"38";
      when x"113" => DATA <= x"66";
      when x"114" => DATA <= x"53";
      when x"115" => DATA <= x"A4";
      when x"116" => DATA <= x"03";
      when x"117" => DATA <= x"88";
      when x"118" => DATA <= x"C8";
      when x"119" => DATA <= x"B1";
      when x"11A" => DATA <= x"05";
      when x"11B" => DATA <= x"C9";
      when x"11C" => DATA <= x"20";
      when x"11D" => DATA <= x"F0";
      when x"11E" => DATA <= x"F9";
      when x"11F" => DATA <= x"88";
      when x"120" => DATA <= x"84";
      when x"121" => DATA <= x"52";
      when x"122" => DATA <= x"CA";
      when x"123" => DATA <= x"A4";
      when x"124" => DATA <= x"52";
      when x"125" => DATA <= x"E8";
      when x"126" => DATA <= x"C8";
      when x"127" => DATA <= x"BD";
      when x"128" => DATA <= x"06";
      when x"129" => DATA <= x"D0";
      when x"12A" => DATA <= x"30";
      when x"12B" => DATA <= x"1A";
      when x"12C" => DATA <= x"D1";
      when x"12D" => DATA <= x"05";
      when x"12E" => DATA <= x"F0";
      when x"12F" => DATA <= x"F5";
      when x"130" => DATA <= x"CA";
      when x"131" => DATA <= x"E8";
      when x"132" => DATA <= x"BD";
      when x"133" => DATA <= x"06";
      when x"134" => DATA <= x"D0";
      when x"135" => DATA <= x"10";
      when x"136" => DATA <= x"FA";
      when x"137" => DATA <= x"E8";
      when x"138" => DATA <= x"24";
      when x"139" => DATA <= x"53";
      when x"13A" => DATA <= x"10";
      when x"13B" => DATA <= x"E7";
      when x"13C" => DATA <= x"B1";
      when x"13D" => DATA <= x"05";
      when x"13E" => DATA <= x"C9";
      when x"13F" => DATA <= x"2E";
      when x"140" => DATA <= x"D0";
      when x"141" => DATA <= x"E1";
      when x"142" => DATA <= x"C8";
      when x"143" => DATA <= x"CA";
      when x"144" => DATA <= x"B0";
      when x"145" => DATA <= x"E1";
      when x"146" => DATA <= x"C9";
      when x"147" => DATA <= x"FE";
      when x"148" => DATA <= x"B0";
      when x"149" => DATA <= x"11";
      when x"14A" => DATA <= x"85";
      when x"14B" => DATA <= x"53";
      when x"14C" => DATA <= x"BD";
      when x"14D" => DATA <= x"07";
      when x"14E" => DATA <= x"D0";
      when x"14F" => DATA <= x"85";
      when x"150" => DATA <= x"52";
      when x"151" => DATA <= x"84";
      when x"152" => DATA <= x"03";
      when x"153" => DATA <= x"A6";
      when x"154" => DATA <= x"04";
      when x"155" => DATA <= x"6C";
      when x"156" => DATA <= x"52";
      when x"157" => DATA <= x"00";
      when x"158" => DATA <= x"A6";
      when x"159" => DATA <= x"04";
      when x"15A" => DATA <= x"60";
      when x"15B" => DATA <= x"F0";
      when x"15C" => DATA <= x"FB";
      when x"15D" => DATA <= x"00";
      when x"15E" => DATA <= x"84";
      when x"15F" => DATA <= x"03";
      when x"160" => DATA <= x"20";
      when x"161" => DATA <= x"EC";
      when x"162" => DATA <= x"D0";
      when x"163" => DATA <= x"20";
      when x"164" => DATA <= x"9A";
      when x"165" => DATA <= x"D8";
      when x"166" => DATA <= x"A5";
      when x"167" => DATA <= x"5A";
      when x"168" => DATA <= x"85";
      when x"169" => DATA <= x"60";
      when x"16A" => DATA <= x"A5";
      when x"16B" => DATA <= x"5B";
      when x"16C" => DATA <= x"85";
      when x"16D" => DATA <= x"5F";
      when x"16E" => DATA <= x"A5";
      when x"16F" => DATA <= x"5C";
      when x"170" => DATA <= x"85";
      when x"171" => DATA <= x"5E";
      when x"172" => DATA <= x"A0";
      when x"173" => DATA <= x"5D";
      when x"174" => DATA <= x"4C";
      when x"175" => DATA <= x"9F";
      when x"176" => DATA <= x"C9";
      when x"177" => DATA <= x"20";
      when x"178" => DATA <= x"F2";
      when x"179" => DATA <= x"D0";
      when x"17A" => DATA <= x"20";
      when x"17B" => DATA <= x"70";
      when x"17C" => DATA <= x"D8";
      when x"17D" => DATA <= x"20";
      when x"17E" => DATA <= x"3C";
      when x"17F" => DATA <= x"D9";
      when x"180" => DATA <= x"4C";
      when x"181" => DATA <= x"FF";
      when x"182" => DATA <= x"D0";
      when x"183" => DATA <= x"20";
      when x"184" => DATA <= x"F2";
      when x"185" => DATA <= x"D0";
      when x"186" => DATA <= x"20";
      when x"187" => DATA <= x"70";
      when x"188" => DATA <= x"D8";
      when x"189" => DATA <= x"20";
      when x"18A" => DATA <= x"39";
      when x"18B" => DATA <= x"D9";
      when x"18C" => DATA <= x"4C";
      when x"18D" => DATA <= x"FF";
      when x"18E" => DATA <= x"D0";
      when x"18F" => DATA <= x"20";
      when x"190" => DATA <= x"03";
      when x"191" => DATA <= x"D1";
      when x"192" => DATA <= x"20";
      when x"193" => DATA <= x"70";
      when x"194" => DATA <= x"D8";
      when x"195" => DATA <= x"20";
      when x"196" => DATA <= x"45";
      when x"197" => DATA <= x"DA";
      when x"198" => DATA <= x"4C";
      when x"199" => DATA <= x"F8";
      when x"19A" => DATA <= x"D0";
      when x"19B" => DATA <= x"20";
      when x"19C" => DATA <= x"03";
      when x"19D" => DATA <= x"D1";
      when x"19E" => DATA <= x"20";
      when x"19F" => DATA <= x"70";
      when x"1A0" => DATA <= x"D8";
      when x"1A1" => DATA <= x"20";
      when x"1A2" => DATA <= x"B6";
      when x"1A3" => DATA <= x"DA";
      when x"1A4" => DATA <= x"4C";
      when x"1A5" => DATA <= x"F8";
      when x"1A6" => DATA <= x"D0";
      when x"1A7" => DATA <= x"20";
      when x"1A8" => DATA <= x"B6";
      when x"1A9" => DATA <= x"DB";
      when x"1AA" => DATA <= x"20";
      when x"1AB" => DATA <= x"5D";
      when x"1AC" => DATA <= x"D8";
      when x"1AD" => DATA <= x"20";
      when x"1AE" => DATA <= x"EB";
      when x"1AF" => DATA <= x"D0";
      when x"1B0" => DATA <= x"20";
      when x"1B1" => DATA <= x"70";
      when x"1B2" => DATA <= x"D8";
      when x"1B3" => DATA <= x"20";
      when x"1B4" => DATA <= x"45";
      when x"1B5" => DATA <= x"DA";
      when x"1B6" => DATA <= x"20";
      when x"1B7" => DATA <= x"D7";
      when x"1B8" => DATA <= x"DD";
      when x"1B9" => DATA <= x"4C";
      when x"1BA" => DATA <= x"09";
      when x"1BB" => DATA <= x"D1";
      when x"1BC" => DATA <= x"20";
      when x"1BD" => DATA <= x"CB";
      when x"1BE" => DATA <= x"D1";
      when x"1BF" => DATA <= x"20";
      when x"1C0" => DATA <= x"86";
      when x"1C1" => DATA <= x"D6";
      when x"1C2" => DATA <= x"F0";
      when x"1C3" => DATA <= x"06";
      when x"1C4" => DATA <= x"A5";
      when x"1C5" => DATA <= x"57";
      when x"1C6" => DATA <= x"49";
      when x"1C7" => DATA <= x"80";
      when x"1C8" => DATA <= x"85";
      when x"1C9" => DATA <= x"57";
      when x"1CA" => DATA <= x"60";
      when x"1CB" => DATA <= x"A4";
      when x"1CC" => DATA <= x"03";
      when x"1CD" => DATA <= x"88";
      when x"1CE" => DATA <= x"C8";
      when x"1CF" => DATA <= x"B1";
      when x"1D0" => DATA <= x"05";
      when x"1D1" => DATA <= x"C9";
      when x"1D2" => DATA <= x"20";
      when x"1D3" => DATA <= x"F0";
      when x"1D4" => DATA <= x"F9";
      when x"1D5" => DATA <= x"C9";
      when x"1D6" => DATA <= x"25";
      when x"1D7" => DATA <= x"D0";
      when x"1D8" => DATA <= x"32";
      when x"1D9" => DATA <= x"E6";
      when x"1DA" => DATA <= x"03";
      when x"1DB" => DATA <= x"20";
      when x"1DC" => DATA <= x"44";
      when x"1DD" => DATA <= x"D4";
      when x"1DE" => DATA <= x"90";
      when x"1DF" => DATA <= x"2B";
      when x"1E0" => DATA <= x"A0";
      when x"1E1" => DATA <= x"6F";
      when x"1E2" => DATA <= x"20";
      when x"1E3" => DATA <= x"CD";
      when x"1E4" => DATA <= x"C3";
      when x"1E5" => DATA <= x"A0";
      when x"1E6" => DATA <= x"04";
      when x"1E7" => DATA <= x"A9";
      when x"1E8" => DATA <= x"00";
      when x"1E9" => DATA <= x"85";
      when x"1EA" => DATA <= x"5E";
      when x"1EB" => DATA <= x"85";
      when x"1EC" => DATA <= x"58";
      when x"1ED" => DATA <= x"85";
      when x"1EE" => DATA <= x"57";
      when x"1EF" => DATA <= x"B1";
      when x"1F0" => DATA <= x"6F";
      when x"1F1" => DATA <= x"99";
      when x"1F2" => DATA <= x"59";
      when x"1F3" => DATA <= x"00";
      when x"1F4" => DATA <= x"05";
      when x"1F5" => DATA <= x"57";
      when x"1F6" => DATA <= x"85";
      when x"1F7" => DATA <= x"57";
      when x"1F8" => DATA <= x"88";
      when x"1F9" => DATA <= x"10";
      when x"1FA" => DATA <= x"F4";
      when x"1FB" => DATA <= x"AA";
      when x"1FC" => DATA <= x"F0";
      when x"1FD" => DATA <= x"09";
      when x"1FE" => DATA <= x"A5";
      when x"1FF" => DATA <= x"5A";
      when x"200" => DATA <= x"85";
      when x"201" => DATA <= x"57";
      when x"202" => DATA <= x"09";
      when x"203" => DATA <= x"80";
      when x"204" => DATA <= x"85";
      when x"205" => DATA <= x"5A";
      when x"206" => DATA <= x"8A";
      when x"207" => DATA <= x"60";
      when x"208" => DATA <= x"84";
      when x"209" => DATA <= x"03";
      when x"20A" => DATA <= x"60";
      when x"20B" => DATA <= x"20";
      when x"20C" => DATA <= x"A5";
      when x"20D" => DATA <= x"D5";
      when x"20E" => DATA <= x"B0";
      when x"20F" => DATA <= x"F8";
      when x"210" => DATA <= x"A2";
      when x"211" => DATA <= x"00";
      when x"212" => DATA <= x"4C";
      when x"213" => DATA <= x"12";
      when x"214" => DATA <= x"D1";
      when x"215" => DATA <= x"20";
      when x"216" => DATA <= x"EB";
      when x"217" => DATA <= x"D0";
      when x"218" => DATA <= x"20";
      when x"219" => DATA <= x"86";
      when x"21A" => DATA <= x"D6";
      when x"21B" => DATA <= x"30";
      when x"21C" => DATA <= x"A7";
      when x"21D" => DATA <= x"60";
      when x"21E" => DATA <= x"20";
      when x"21F" => DATA <= x"24";
      when x"220" => DATA <= x"D2";
      when x"221" => DATA <= x"4C";
      when x"222" => DATA <= x"86";
      when x"223" => DATA <= x"DC";
      when x"224" => DATA <= x"20";
      when x"225" => DATA <= x"EB";
      when x"226" => DATA <= x"D0";
      when x"227" => DATA <= x"20";
      when x"228" => DATA <= x"86";
      when x"229" => DATA <= x"D6";
      when x"22A" => DATA <= x"10";
      when x"22B" => DATA <= x"0A";
      when x"22C" => DATA <= x"A9";
      when x"22D" => DATA <= x"00";
      when x"22E" => DATA <= x"85";
      when x"22F" => DATA <= x"57";
      when x"230" => DATA <= x"20";
      when x"231" => DATA <= x"36";
      when x"232" => DATA <= x"D2";
      when x"233" => DATA <= x"4C";
      when x"234" => DATA <= x"75";
      when x"235" => DATA <= x"DC";
      when x"236" => DATA <= x"20";
      when x"237" => DATA <= x"2C";
      when x"238" => DATA <= x"D8";
      when x"239" => DATA <= x"20";
      when x"23A" => DATA <= x"45";
      when x"23B" => DATA <= x"DA";
      when x"23C" => DATA <= x"20";
      when x"23D" => DATA <= x"31";
      when x"23E" => DATA <= x"D8";
      when x"23F" => DATA <= x"20";
      when x"240" => DATA <= x"8D";
      when x"241" => DATA <= x"DE";
      when x"242" => DATA <= x"20";
      when x"243" => DATA <= x"33";
      when x"244" => DATA <= x"D9";
      when x"245" => DATA <= x"20";
      when x"246" => DATA <= x"72";
      when x"247" => DATA <= x"DB";
      when x"248" => DATA <= x"20";
      when x"249" => DATA <= x"86";
      when x"24A" => DATA <= x"D6";
      when x"24B" => DATA <= x"F0";
      when x"24C" => DATA <= x"12";
      when x"24D" => DATA <= x"20";
      when x"24E" => DATA <= x"31";
      when x"24F" => DATA <= x"D8";
      when x"250" => DATA <= x"20";
      when x"251" => DATA <= x"A6";
      when x"252" => DATA <= x"DB";
      when x"253" => DATA <= x"20";
      when x"254" => DATA <= x"E5";
      when x"255" => DATA <= x"D1";
      when x"256" => DATA <= x"20";
      when x"257" => DATA <= x"AA";
      when x"258" => DATA <= x"DB";
      when x"259" => DATA <= x"20";
      when x"25A" => DATA <= x"DC";
      when x"25B" => DATA <= x"DA";
      when x"25C" => DATA <= x"4C";
      when x"25D" => DATA <= x"67";
      when x"25E" => DATA <= x"DC";
      when x"25F" => DATA <= x"20";
      when x"260" => DATA <= x"93";
      when x"261" => DATA <= x"DD";
      when x"262" => DATA <= x"4C";
      when x"263" => DATA <= x"E5";
      when x"264" => DATA <= x"D1";
      when x"265" => DATA <= x"20";
      when x"266" => DATA <= x"EB";
      when x"267" => DATA <= x"D0";
      when x"268" => DATA <= x"A0";
      when x"269" => DATA <= x"7C";
      when x"26A" => DATA <= x"A9";
      when x"26B" => DATA <= x"D2";
      when x"26C" => DATA <= x"84";
      when x"26D" => DATA <= x"6F";
      when x"26E" => DATA <= x"85";
      when x"26F" => DATA <= x"70";
      when x"270" => DATA <= x"4C";
      when x"271" => DATA <= x"45";
      when x"272" => DATA <= x"DA";
      when x"273" => DATA <= x"20";
      when x"274" => DATA <= x"EB";
      when x"275" => DATA <= x"D0";
      when x"276" => DATA <= x"A0";
      when x"277" => DATA <= x"81";
      when x"278" => DATA <= x"A9";
      when x"279" => DATA <= x"D2";
      when x"27A" => DATA <= x"D0";
      when x"27B" => DATA <= x"F0";
      when x"27C" => DATA <= x"7B";
      when x"27D" => DATA <= x"0E";
      when x"27E" => DATA <= x"FA";
      when x"27F" => DATA <= x"35";
      when x"280" => DATA <= x"12";
      when x"281" => DATA <= x"86";
      when x"282" => DATA <= x"65";
      when x"283" => DATA <= x"2E";
      when x"284" => DATA <= x"E0";
      when x"285" => DATA <= x"D3";
      when x"286" => DATA <= x"20";
      when x"287" => DATA <= x"EB";
      when x"288" => DATA <= x"D0";
      when x"289" => DATA <= x"20";
      when x"28A" => DATA <= x"86";
      when x"28B" => DATA <= x"D6";
      when x"28C" => DATA <= x"F0";
      when x"28D" => DATA <= x"07";
      when x"28E" => DATA <= x"48";
      when x"28F" => DATA <= x"20";
      when x"290" => DATA <= x"8D";
      when x"291" => DATA <= x"DE";
      when x"292" => DATA <= x"68";
      when x"293" => DATA <= x"85";
      when x"294" => DATA <= x"57";
      when x"295" => DATA <= x"60";
      when x"296" => DATA <= x"24";
      when x"297" => DATA <= x"73";
      when x"298" => DATA <= x"30";
      when x"299" => DATA <= x"26";
      when x"29A" => DATA <= x"20";
      when x"29B" => DATA <= x"BC";
      when x"29C" => DATA <= x"C8";
      when x"29D" => DATA <= x"A0";
      when x"29E" => DATA <= x"5D";
      when x"29F" => DATA <= x"20";
      when x"2A0" => DATA <= x"CD";
      when x"2A1" => DATA <= x"C3";
      when x"2A2" => DATA <= x"85";
      when x"2A3" => DATA <= x"5A";
      when x"2A4" => DATA <= x"A5";
      when x"2A5" => DATA <= x"5F";
      when x"2A6" => DATA <= x"85";
      when x"2A7" => DATA <= x"5B";
      when x"2A8" => DATA <= x"A5";
      when x"2A9" => DATA <= x"5E";
      when x"2AA" => DATA <= x"85";
      when x"2AB" => DATA <= x"5C";
      when x"2AC" => DATA <= x"A9";
      when x"2AD" => DATA <= x"A0";
      when x"2AE" => DATA <= x"85";
      when x"2AF" => DATA <= x"59";
      when x"2B0" => DATA <= x"A0";
      when x"2B1" => DATA <= x"00";
      when x"2B2" => DATA <= x"84";
      when x"2B3" => DATA <= x"5E";
      when x"2B4" => DATA <= x"A5";
      when x"2B5" => DATA <= x"5A";
      when x"2B6" => DATA <= x"85";
      when x"2B7" => DATA <= x"57";
      when x"2B8" => DATA <= x"10";
      when x"2B9" => DATA <= x"03";
      when x"2BA" => DATA <= x"20";
      when x"2BB" => DATA <= x"D5";
      when x"2BC" => DATA <= x"D8";
      when x"2BD" => DATA <= x"4C";
      when x"2BE" => DATA <= x"C8";
      when x"2BF" => DATA <= x"D7";
      when x"2C0" => DATA <= x"4C";
      when x"2C1" => DATA <= x"1B";
      when x"2C2" => DATA <= x"CA";
      when x"2C3" => DATA <= x"20";
      when x"2C4" => DATA <= x"93";
      when x"2C5" => DATA <= x"DD";
      when x"2C6" => DATA <= x"20";
      when x"2C7" => DATA <= x"E5";
      when x"2C8" => DATA <= x"D1";
      when x"2C9" => DATA <= x"E6";
      when x"2CA" => DATA <= x"59";
      when x"2CB" => DATA <= x"60";
      when x"2CC" => DATA <= x"20";
      when x"2CD" => DATA <= x"3E";
      when x"2CE" => DATA <= x"CF";
      when x"2CF" => DATA <= x"A2";
      when x"2D0" => DATA <= x"04";
      when x"2D1" => DATA <= x"20";
      when x"2D2" => DATA <= x"D4";
      when x"2D3" => DATA <= x"FF";
      when x"2D4" => DATA <= x"9D";
      when x"2D5" => DATA <= x"C5";
      when x"2D6" => DATA <= x"03";
      when x"2D7" => DATA <= x"CA";
      when x"2D8" => DATA <= x"10";
      when x"2D9" => DATA <= x"F7";
      when x"2DA" => DATA <= x"20";
      when x"2DB" => DATA <= x"AA";
      when x"2DC" => DATA <= x"DB";
      when x"2DD" => DATA <= x"4C";
      when x"2DE" => DATA <= x"E5";
      when x"2DF" => DATA <= x"D1";
      when x"2E0" => DATA <= x"20";
      when x"2E1" => DATA <= x"B1";
      when x"2E2" => DATA <= x"CE";
      when x"2E3" => DATA <= x"A0";
      when x"2E4" => DATA <= x"00";
      when x"2E5" => DATA <= x"20";
      when x"2E6" => DATA <= x"04";
      when x"2E7" => DATA <= x"D3";
      when x"2E8" => DATA <= x"C9";
      when x"2E9" => DATA <= x"2B";
      when x"2EA" => DATA <= x"F0";
      when x"2EB" => DATA <= x"0F";
      when x"2EC" => DATA <= x"C9";
      when x"2ED" => DATA <= x"2D";
      when x"2EE" => DATA <= x"D0";
      when x"2EF" => DATA <= x"0E";
      when x"2F0" => DATA <= x"20";
      when x"2F1" => DATA <= x"03";
      when x"2F2" => DATA <= x"D3";
      when x"2F3" => DATA <= x"84";
      when x"2F4" => DATA <= x"54";
      when x"2F5" => DATA <= x"20";
      when x"2F6" => DATA <= x"B1";
      when x"2F7" => DATA <= x"D5";
      when x"2F8" => DATA <= x"4C";
      when x"2F9" => DATA <= x"BF";
      when x"2FA" => DATA <= x"D1";
      when x"2FB" => DATA <= x"20";
      when x"2FC" => DATA <= x"03";
      when x"2FD" => DATA <= x"D3";
      when x"2FE" => DATA <= x"84";
      when x"2FF" => DATA <= x"54";
      when x"300" => DATA <= x"4C";
      when x"301" => DATA <= x"B1";
      when x"302" => DATA <= x"D5";
      when x"303" => DATA <= x"C8";
      when x"304" => DATA <= x"B1";
      when x"305" => DATA <= x"52";
      when x"306" => DATA <= x"C9";
      when x"307" => DATA <= x"20";
      when x"308" => DATA <= x"F0";
      when x"309" => DATA <= x"F9";
      when x"30A" => DATA <= x"60";
      when x"30B" => DATA <= x"20";
      when x"30C" => DATA <= x"44";
      when x"30D" => DATA <= x"D4";
      when x"30E" => DATA <= x"90";
      when x"30F" => DATA <= x"D4";
      when x"310" => DATA <= x"20";
      when x"311" => DATA <= x"79";
      when x"312" => DATA <= x"C2";
      when x"313" => DATA <= x"20";
      when x"314" => DATA <= x"FC";
      when x"315" => DATA <= x"D0";
      when x"316" => DATA <= x"20";
      when x"317" => DATA <= x"E4";
      when x"318" => DATA <= x"C4";
      when x"319" => DATA <= x"20";
      when x"31A" => DATA <= x"36";
      when x"31B" => DATA <= x"D8";
      when x"31C" => DATA <= x"4C";
      when x"31D" => DATA <= x"5B";
      when x"31E" => DATA <= x"C5";
      when x"31F" => DATA <= x"20";
      when x"320" => DATA <= x"FC";
      when x"321" => DATA <= x"D0";
      when x"322" => DATA <= x"20";
      when x"323" => DATA <= x"31";
      when x"324" => DATA <= x"C2";
      when x"325" => DATA <= x"20";
      when x"326" => DATA <= x"E1";
      when x"327" => DATA <= x"C4";
      when x"328" => DATA <= x"20";
      when x"329" => DATA <= x"CB";
      when x"32A" => DATA <= x"C3";
      when x"32B" => DATA <= x"20";
      when x"32C" => DATA <= x"D0";
      when x"32D" => DATA <= x"D4";
      when x"32E" => DATA <= x"4C";
      when x"32F" => DATA <= x"5B";
      when x"330" => DATA <= x"C5";
      when x"331" => DATA <= x"20";
      when x"332" => DATA <= x"72";
      when x"333" => DATA <= x"C3";
      when x"334" => DATA <= x"A2";
      when x"335" => DATA <= x"B8";
      when x"336" => DATA <= x"4C";
      when x"337" => DATA <= x"0B";
      when x"338" => DATA <= x"D1";
      when x"339" => DATA <= x"20";
      when x"33A" => DATA <= x"FC";
      when x"33B" => DATA <= x"D0";
      when x"33C" => DATA <= x"A9";
      when x"33D" => DATA <= x"C5";
      when x"33E" => DATA <= x"85";
      when x"33F" => DATA <= x"52";
      when x"340" => DATA <= x"A9";
      when x"341" => DATA <= x"03";
      when x"342" => DATA <= x"85";
      when x"343" => DATA <= x"53";
      when x"344" => DATA <= x"20";
      when x"345" => DATA <= x"D0";
      when x"346" => DATA <= x"D4";
      when x"347" => DATA <= x"C6";
      when x"348" => DATA <= x"6F";
      when x"349" => DATA <= x"AD";
      when x"34A" => DATA <= x"21";
      when x"34B" => DATA <= x"03";
      when x"34C" => DATA <= x"38";
      when x"34D" => DATA <= x"E5";
      when x"34E" => DATA <= x"6F";
      when x"34F" => DATA <= x"90";
      when x"350" => DATA <= x"0B";
      when x"351" => DATA <= x"F0";
      when x"352" => DATA <= x"09";
      when x"353" => DATA <= x"A8";
      when x"354" => DATA <= x"A9";
      when x"355" => DATA <= x"20";
      when x"356" => DATA <= x"20";
      when x"357" => DATA <= x"4C";
      when x"358" => DATA <= x"CA";
      when x"359" => DATA <= x"88";
      when x"35A" => DATA <= x"D0";
      when x"35B" => DATA <= x"FA";
      when x"35C" => DATA <= x"A0";
      when x"35D" => DATA <= x"00";
      when x"35E" => DATA <= x"B1";
      when x"35F" => DATA <= x"52";
      when x"360" => DATA <= x"C9";
      when x"361" => DATA <= x"0D";
      when x"362" => DATA <= x"F0";
      when x"363" => DATA <= x"CD";
      when x"364" => DATA <= x"20";
      when x"365" => DATA <= x"4C";
      when x"366" => DATA <= x"CA";
      when x"367" => DATA <= x"C8";
      when x"368" => DATA <= x"D0";
      when x"369" => DATA <= x"F4";
      when x"36A" => DATA <= x"20";
      when x"36B" => DATA <= x"72";
      when x"36C" => DATA <= x"C3";
      when x"36D" => DATA <= x"B1";
      when x"36E" => DATA <= x"05";
      when x"36F" => DATA <= x"C9";
      when x"370" => DATA <= x"25";
      when x"371" => DATA <= x"D0";
      when x"372" => DATA <= x"08";
      when x"373" => DATA <= x"C8";
      when x"374" => DATA <= x"84";
      when x"375" => DATA <= x"03";
      when x"376" => DATA <= x"20";
      when x"377" => DATA <= x"44";
      when x"378" => DATA <= x"D4";
      when x"379" => DATA <= x"B0";
      when x"37A" => DATA <= x"05";
      when x"37B" => DATA <= x"A2";
      when x"37C" => DATA <= x"C3";
      when x"37D" => DATA <= x"4C";
      when x"37E" => DATA <= x"0B";
      when x"37F" => DATA <= x"D1";
      when x"380" => DATA <= x"20";
      when x"381" => DATA <= x"09";
      when x"382" => DATA <= x"CD";
      when x"383" => DATA <= x"A8";
      when x"384" => DATA <= x"A5";
      when x"385" => DATA <= x"05";
      when x"386" => DATA <= x"48";
      when x"387" => DATA <= x"A5";
      when x"388" => DATA <= x"06";
      when x"389" => DATA <= x"48";
      when x"38A" => DATA <= x"A5";
      when x"38B" => DATA <= x"03";
      when x"38C" => DATA <= x"48";
      when x"38D" => DATA <= x"84";
      when x"38E" => DATA <= x"03";
      when x"38F" => DATA <= x"C8";
      when x"390" => DATA <= x"84";
      when x"391" => DATA <= x"06";
      when x"392" => DATA <= x"A9";
      when x"393" => DATA <= x"40";
      when x"394" => DATA <= x"85";
      when x"395" => DATA <= x"05";
      when x"396" => DATA <= x"20";
      when x"397" => DATA <= x"FC";
      when x"398" => DATA <= x"D0";
      when x"399" => DATA <= x"68";
      when x"39A" => DATA <= x"85";
      when x"39B" => DATA <= x"03";
      when x"39C" => DATA <= x"68";
      when x"39D" => DATA <= x"85";
      when x"39E" => DATA <= x"06";
      when x"39F" => DATA <= x"68";
      when x"3A0" => DATA <= x"85";
      when x"3A1" => DATA <= x"05";
      when x"3A2" => DATA <= x"20";
      when x"3A3" => DATA <= x"36";
      when x"3A4" => DATA <= x"D8";
      when x"3A5" => DATA <= x"4C";
      when x"3A6" => DATA <= x"7B";
      when x"3A7" => DATA <= x"D3";
      when x"3A8" => DATA <= x"20";
      when x"3A9" => DATA <= x"EB";
      when x"3AA" => DATA <= x"D9";
      when x"3AB" => DATA <= x"4C";
      when x"3AC" => DATA <= x"69";
      when x"3AD" => DATA <= x"C5";
      when x"3AE" => DATA <= x"20";
      when x"3AF" => DATA <= x"EB";
      when x"3B0" => DATA <= x"D9";
      when x"3B1" => DATA <= x"4C";
      when x"3B2" => DATA <= x"D5";
      when x"3B3" => DATA <= x"CC";
      when x"3B4" => DATA <= x"20";
      when x"3B5" => DATA <= x"94";
      when x"3B6" => DATA <= x"D4";
      when x"3B7" => DATA <= x"20";
      when x"3B8" => DATA <= x"FC";
      when x"3B9" => DATA <= x"D0";
      when x"3BA" => DATA <= x"20";
      when x"3BB" => DATA <= x"E4";
      when x"3BC" => DATA <= x"C4";
      when x"3BD" => DATA <= x"20";
      when x"3BE" => DATA <= x"31";
      when x"3BF" => DATA <= x"D8";
      when x"3C0" => DATA <= x"A6";
      when x"3C1" => DATA <= x"04";
      when x"3C2" => DATA <= x"20";
      when x"3C3" => DATA <= x"41";
      when x"3C4" => DATA <= x"CF";
      when x"3C5" => DATA <= x"A2";
      when x"3C6" => DATA <= x"04";
      when x"3C7" => DATA <= x"BD";
      when x"3C8" => DATA <= x"C5";
      when x"3C9" => DATA <= x"03";
      when x"3CA" => DATA <= x"20";
      when x"3CB" => DATA <= x"D1";
      when x"3CC" => DATA <= x"FF";
      when x"3CD" => DATA <= x"CA";
      when x"3CE" => DATA <= x"10";
      when x"3CF" => DATA <= x"F7";
      when x"3D0" => DATA <= x"4C";
      when x"3D1" => DATA <= x"5B";
      when x"3D2" => DATA <= x"C5";
      when x"3D3" => DATA <= x"A5";
      when x"3D4" => DATA <= x"01";
      when x"3D5" => DATA <= x"05";
      when x"3D6" => DATA <= x"02";
      when x"3D7" => DATA <= x"F0";
      when x"3D8" => DATA <= x"6A";
      when x"3D9" => DATA <= x"20";
      when x"3DA" => DATA <= x"34";
      when x"3DB" => DATA <= x"C4";
      when x"3DC" => DATA <= x"B0";
      when x"3DD" => DATA <= x"65";
      when x"3DE" => DATA <= x"A4";
      when x"3DF" => DATA <= x"03";
      when x"3E0" => DATA <= x"B1";
      when x"3E1" => DATA <= x"05";
      when x"3E2" => DATA <= x"C9";
      when x"3E3" => DATA <= x"25";
      when x"3E4" => DATA <= x"D0";
      when x"3E5" => DATA <= x"5D";
      when x"3E6" => DATA <= x"C8";
      when x"3E7" => DATA <= x"B1";
      when x"3E8" => DATA <= x"05";
      when x"3E9" => DATA <= x"C8";
      when x"3EA" => DATA <= x"D1";
      when x"3EB" => DATA <= x"05";
      when x"3EC" => DATA <= x"D0";
      when x"3ED" => DATA <= x"55";
      when x"3EE" => DATA <= x"C9";
      when x"3EF" => DATA <= x"5B";
      when x"3F0" => DATA <= x"B0";
      when x"3F1" => DATA <= x"51";
      when x"3F2" => DATA <= x"E9";
      when x"3F3" => DATA <= x"3F";
      when x"3F4" => DATA <= x"90";
      when x"3F5" => DATA <= x"4D";
      when x"3F6" => DATA <= x"C8";
      when x"3F7" => DATA <= x"84";
      when x"3F8" => DATA <= x"03";
      when x"3F9" => DATA <= x"48";
      when x"3FA" => DATA <= x"20";
      when x"3FB" => DATA <= x"8B";
      when x"3FC" => DATA <= x"C7";
      when x"3FD" => DATA <= x"F6";
      when x"3FE" => DATA <= x"15";
      when x"3FF" => DATA <= x"D0";
      when x"400" => DATA <= x"02";
      when x"401" => DATA <= x"F6";
      when x"402" => DATA <= x"24";
      when x"403" => DATA <= x"20";
      when x"404" => DATA <= x"9A";
      when x"405" => DATA <= x"D4";
      when x"406" => DATA <= x"68";
      when x"407" => DATA <= x"A8";
      when x"408" => DATA <= x"18";
      when x"409" => DATA <= x"A5";
      when x"40A" => DATA <= x"23";
      when x"40B" => DATA <= x"99";
      when x"40C" => DATA <= x"87";
      when x"40D" => DATA <= x"28";
      when x"40E" => DATA <= x"65";
      when x"40F" => DATA <= x"16";
      when x"410" => DATA <= x"85";
      when x"411" => DATA <= x"23";
      when x"412" => DATA <= x"A5";
      when x"413" => DATA <= x"24";
      when x"414" => DATA <= x"99";
      when x"415" => DATA <= x"A2";
      when x"416" => DATA <= x"28";
      when x"417" => DATA <= x"65";
      when x"418" => DATA <= x"25";
      when x"419" => DATA <= x"85";
      when x"41A" => DATA <= x"24";
      when x"41B" => DATA <= x"A0";
      when x"41C" => DATA <= x"00";
      when x"41D" => DATA <= x"84";
      when x"41E" => DATA <= x"04";
      when x"41F" => DATA <= x"A9";
      when x"420" => DATA <= x"AA";
      when x"421" => DATA <= x"91";
      when x"422" => DATA <= x"23";
      when x"423" => DATA <= x"D1";
      when x"424" => DATA <= x"23";
      when x"425" => DATA <= x"D0";
      when x"426" => DATA <= x"1C";
      when x"427" => DATA <= x"4A";
      when x"428" => DATA <= x"91";
      when x"429" => DATA <= x"23";
      when x"42A" => DATA <= x"D1";
      when x"42B" => DATA <= x"23";
      when x"42C" => DATA <= x"D0";
      when x"42D" => DATA <= x"15";
      when x"42E" => DATA <= x"20";
      when x"42F" => DATA <= x"34";
      when x"430" => DATA <= x"C4";
      when x"431" => DATA <= x"B0";
      when x"432" => DATA <= x"10";
      when x"433" => DATA <= x"A4";
      when x"434" => DATA <= x"03";
      when x"435" => DATA <= x"B1";
      when x"436" => DATA <= x"05";
      when x"437" => DATA <= x"C9";
      when x"438" => DATA <= x"2C";
      when x"439" => DATA <= x"D0";
      when x"43A" => DATA <= x"05";
      when x"43B" => DATA <= x"E6";
      when x"43C" => DATA <= x"03";
      when x"43D" => DATA <= x"4C";
      when x"43E" => DATA <= x"D3";
      when x"43F" => DATA <= x"D3";
      when x"440" => DATA <= x"4C";
      when x"441" => DATA <= x"58";
      when x"442" => DATA <= x"C5";
      when x"443" => DATA <= x"00";
      when x"444" => DATA <= x"20";
      when x"445" => DATA <= x"34";
      when x"446" => DATA <= x"C4";
      when x"447" => DATA <= x"90";
      when x"448" => DATA <= x"0E";
      when x"449" => DATA <= x"B5";
      when x"44A" => DATA <= x"15";
      when x"44B" => DATA <= x"0A";
      when x"44C" => DATA <= x"0A";
      when x"44D" => DATA <= x"75";
      when x"44E" => DATA <= x"15";
      when x"44F" => DATA <= x"95";
      when x"450" => DATA <= x"15";
      when x"451" => DATA <= x"A9";
      when x"452" => DATA <= x"28";
      when x"453" => DATA <= x"95";
      when x"454" => DATA <= x"24";
      when x"455" => DATA <= x"38";
      when x"456" => DATA <= x"60";
      when x"457" => DATA <= x"A4";
      when x"458" => DATA <= x"03";
      when x"459" => DATA <= x"B1";
      when x"45A" => DATA <= x"05";
      when x"45B" => DATA <= x"C9";
      when x"45C" => DATA <= x"21";
      when x"45D" => DATA <= x"D0";
      when x"45E" => DATA <= x"07";
      when x"45F" => DATA <= x"E6";
      when x"460" => DATA <= x"03";
      when x"461" => DATA <= x"20";
      when x"462" => DATA <= x"BC";
      when x"463" => DATA <= x"C8";
      when x"464" => DATA <= x"38";
      when x"465" => DATA <= x"60";
      when x"466" => DATA <= x"C8";
      when x"467" => DATA <= x"D1";
      when x"468" => DATA <= x"05";
      when x"469" => DATA <= x"D0";
      when x"46A" => DATA <= x"08";
      when x"46B" => DATA <= x"C9";
      when x"46C" => DATA <= x"5B";
      when x"46D" => DATA <= x"B0";
      when x"46E" => DATA <= x"04";
      when x"46F" => DATA <= x"E9";
      when x"470" => DATA <= x"3F";
      when x"471" => DATA <= x"B0";
      when x"472" => DATA <= x"02";
      when x"473" => DATA <= x"18";
      when x"474" => DATA <= x"60";
      when x"475" => DATA <= x"C8";
      when x"476" => DATA <= x"84";
      when x"477" => DATA <= x"03";
      when x"478" => DATA <= x"48";
      when x"479" => DATA <= x"20";
      when x"47A" => DATA <= x"BC";
      when x"47B" => DATA <= x"C8";
      when x"47C" => DATA <= x"20";
      when x"47D" => DATA <= x"9A";
      when x"47E" => DATA <= x"D4";
      when x"47F" => DATA <= x"68";
      when x"480" => DATA <= x"A8";
      when x"481" => DATA <= x"B0";
      when x"482" => DATA <= x"10";
      when x"483" => DATA <= x"B9";
      when x"484" => DATA <= x"87";
      when x"485" => DATA <= x"28";
      when x"486" => DATA <= x"75";
      when x"487" => DATA <= x"15";
      when x"488" => DATA <= x"95";
      when x"489" => DATA <= x"15";
      when x"48A" => DATA <= x"B9";
      when x"48B" => DATA <= x"A2";
      when x"48C" => DATA <= x"28";
      when x"48D" => DATA <= x"75";
      when x"48E" => DATA <= x"24";
      when x"48F" => DATA <= x"95";
      when x"490" => DATA <= x"24";
      when x"491" => DATA <= x"90";
      when x"492" => DATA <= x"D1";
      when x"493" => DATA <= x"00";
      when x"494" => DATA <= x"20";
      when x"495" => DATA <= x"BC";
      when x"496" => DATA <= x"C8";
      when x"497" => DATA <= x"4C";
      when x"498" => DATA <= x"31";
      when x"499" => DATA <= x"C2";
      when x"49A" => DATA <= x"B4";
      when x"49B" => DATA <= x"24";
      when x"49C" => DATA <= x"B5";
      when x"49D" => DATA <= x"15";
      when x"49E" => DATA <= x"0A";
      when x"49F" => DATA <= x"36";
      when x"4A0" => DATA <= x"24";
      when x"4A1" => DATA <= x"0A";
      when x"4A2" => DATA <= x"36";
      when x"4A3" => DATA <= x"24";
      when x"4A4" => DATA <= x"18";
      when x"4A5" => DATA <= x"75";
      when x"4A6" => DATA <= x"15";
      when x"4A7" => DATA <= x"95";
      when x"4A8" => DATA <= x"15";
      when x"4A9" => DATA <= x"98";
      when x"4AA" => DATA <= x"75";
      when x"4AB" => DATA <= x"24";
      when x"4AC" => DATA <= x"95";
      when x"4AD" => DATA <= x"24";
      when x"4AE" => DATA <= x"60";
      when x"4AF" => DATA <= x"AD";
      when x"4B0" => DATA <= x"04";
      when x"4B1" => DATA <= x"E0";
      when x"4B2" => DATA <= x"C9";
      when x"4B3" => DATA <= x"BF";
      when x"4B4" => DATA <= x"F0";
      when x"4B5" => DATA <= x"0A";
      when x"4B6" => DATA <= x"AD";
      when x"4B7" => DATA <= x"00";
      when x"4B8" => DATA <= x"A0";
      when x"4B9" => DATA <= x"C9";
      when x"4BA" => DATA <= x"40";
      when x"4BB" => DATA <= x"D0";
      when x"4BC" => DATA <= x"83";
      when x"4BD" => DATA <= x"4C";
      when x"4BE" => DATA <= x"02";
      when x"4BF" => DATA <= x"A0";
      when x"4C0" => DATA <= x"4C";
      when x"4C1" => DATA <= x"05";
      when x"4C2" => DATA <= x"E0";
      when x"4C3" => DATA <= x"C9";
      when x"4C4" => DATA <= x"3A";
      when x"4C5" => DATA <= x"B0";
      when x"4C6" => DATA <= x"07";
      when x"4C7" => DATA <= x"C9";
      when x"4C8" => DATA <= x"30";
      when x"4C9" => DATA <= x"90";
      when x"4CA" => DATA <= x"02";
      when x"4CB" => DATA <= x"E9";
      when x"4CC" => DATA <= x"30";
      when x"4CD" => DATA <= x"60";
      when x"4CE" => DATA <= x"18";
      when x"4CF" => DATA <= x"60";
      when x"4D0" => DATA <= x"A9";
      when x"4D1" => DATA <= x"00";
      when x"4D2" => DATA <= x"85";
      when x"4D3" => DATA <= x"6F";
      when x"4D4" => DATA <= x"20";
      when x"4D5" => DATA <= x"86";
      when x"4D6" => DATA <= x"D6";
      when x"4D7" => DATA <= x"D0";
      when x"4D8" => DATA <= x"12";
      when x"4D9" => DATA <= x"A9";
      when x"4DA" => DATA <= x"30";
      when x"4DB" => DATA <= x"20";
      when x"4DC" => DATA <= x"8D";
      when x"4DD" => DATA <= x"D5";
      when x"4DE" => DATA <= x"A9";
      when x"4DF" => DATA <= x"2E";
      when x"4E0" => DATA <= x"20";
      when x"4E1" => DATA <= x"8D";
      when x"4E2" => DATA <= x"D5";
      when x"4E3" => DATA <= x"A9";
      when x"4E4" => DATA <= x"30";
      when x"4E5" => DATA <= x"20";
      when x"4E6" => DATA <= x"8D";
      when x"4E7" => DATA <= x"D5";
      when x"4E8" => DATA <= x"4C";
      when x"4E9" => DATA <= x"71";
      when x"4EA" => DATA <= x"D5";
      when x"4EB" => DATA <= x"10";
      when x"4EC" => DATA <= x"05";
      when x"4ED" => DATA <= x"A9";
      when x"4EE" => DATA <= x"2D";
      when x"4EF" => DATA <= x"20";
      when x"4F0" => DATA <= x"8D";
      when x"4F1" => DATA <= x"D5";
      when x"4F2" => DATA <= x"A9";
      when x"4F3" => DATA <= x"00";
      when x"4F4" => DATA <= x"85";
      when x"4F5" => DATA <= x"6D";
      when x"4F6" => DATA <= x"A5";
      when x"4F7" => DATA <= x"59";
      when x"4F8" => DATA <= x"C9";
      when x"4F9" => DATA <= x"81";
      when x"4FA" => DATA <= x"B0";
      when x"4FB" => DATA <= x"08";
      when x"4FC" => DATA <= x"20";
      when x"4FD" => DATA <= x"A0";
      when x"4FE" => DATA <= x"D6";
      when x"4FF" => DATA <= x"C6";
      when x"500" => DATA <= x"6D";
      when x"501" => DATA <= x"4C";
      when x"502" => DATA <= x"F6";
      when x"503" => DATA <= x"D4";
      when x"504" => DATA <= x"C9";
      when x"505" => DATA <= x"84";
      when x"506" => DATA <= x"90";
      when x"507" => DATA <= x"10";
      when x"508" => DATA <= x"D0";
      when x"509" => DATA <= x"06";
      when x"50A" => DATA <= x"A5";
      when x"50B" => DATA <= x"5A";
      when x"50C" => DATA <= x"C9";
      when x"50D" => DATA <= x"A0";
      when x"50E" => DATA <= x"90";
      when x"50F" => DATA <= x"08";
      when x"510" => DATA <= x"20";
      when x"511" => DATA <= x"1B";
      when x"512" => DATA <= x"D7";
      when x"513" => DATA <= x"E6";
      when x"514" => DATA <= x"6D";
      when x"515" => DATA <= x"4C";
      when x"516" => DATA <= x"F6";
      when x"517" => DATA <= x"D4";
      when x"518" => DATA <= x"A5";
      when x"519" => DATA <= x"59";
      when x"51A" => DATA <= x"C9";
      when x"51B" => DATA <= x"84";
      when x"51C" => DATA <= x"B0";
      when x"51D" => DATA <= x"07";
      when x"51E" => DATA <= x"20";
      when x"51F" => DATA <= x"D8";
      when x"520" => DATA <= x"D6";
      when x"521" => DATA <= x"E6";
      when x"522" => DATA <= x"59";
      when x"523" => DATA <= x"D0";
      when x"524" => DATA <= x"F3";
      when x"525" => DATA <= x"38";
      when x"526" => DATA <= x"A9";
      when x"527" => DATA <= x"FF";
      when x"528" => DATA <= x"20";
      when x"529" => DATA <= x"36";
      when x"52A" => DATA <= x"D6";
      when x"52B" => DATA <= x"A5";
      when x"52C" => DATA <= x"5A";
      when x"52D" => DATA <= x"C9";
      when x"52E" => DATA <= x"A0";
      when x"52F" => DATA <= x"B0";
      when x"530" => DATA <= x"DF";
      when x"531" => DATA <= x"A9";
      when x"532" => DATA <= x"01";
      when x"533" => DATA <= x"A4";
      when x"534" => DATA <= x"6D";
      when x"535" => DATA <= x"30";
      when x"536" => DATA <= x"0A";
      when x"537" => DATA <= x"C0";
      when x"538" => DATA <= x"08";
      when x"539" => DATA <= x"B0";
      when x"53A" => DATA <= x"06";
      when x"53B" => DATA <= x"C8";
      when x"53C" => DATA <= x"A9";
      when x"53D" => DATA <= x"00";
      when x"53E" => DATA <= x"85";
      when x"53F" => DATA <= x"6D";
      when x"540" => DATA <= x"98";
      when x"541" => DATA <= x"85";
      when x"542" => DATA <= x"70";
      when x"543" => DATA <= x"A2";
      when x"544" => DATA <= x"09";
      when x"545" => DATA <= x"86";
      when x"546" => DATA <= x"54";
      when x"547" => DATA <= x"20";
      when x"548" => DATA <= x"75";
      when x"549" => DATA <= x"D5";
      when x"54A" => DATA <= x"C6";
      when x"54B" => DATA <= x"70";
      when x"54C" => DATA <= x"D0";
      when x"54D" => DATA <= x"05";
      when x"54E" => DATA <= x"A9";
      when x"54F" => DATA <= x"2E";
      when x"550" => DATA <= x"20";
      when x"551" => DATA <= x"8D";
      when x"552" => DATA <= x"D5";
      when x"553" => DATA <= x"C6";
      when x"554" => DATA <= x"54";
      when x"555" => DATA <= x"D0";
      when x"556" => DATA <= x"F0";
      when x"557" => DATA <= x"A5";
      when x"558" => DATA <= x"6D";
      when x"559" => DATA <= x"F0";
      when x"55A" => DATA <= x"16";
      when x"55B" => DATA <= x"A9";
      when x"55C" => DATA <= x"45";
      when x"55D" => DATA <= x"20";
      when x"55E" => DATA <= x"8D";
      when x"55F" => DATA <= x"D5";
      when x"560" => DATA <= x"A5";
      when x"561" => DATA <= x"6D";
      when x"562" => DATA <= x"10";
      when x"563" => DATA <= x"0A";
      when x"564" => DATA <= x"A9";
      when x"565" => DATA <= x"2D";
      when x"566" => DATA <= x"20";
      when x"567" => DATA <= x"8D";
      when x"568" => DATA <= x"D5";
      when x"569" => DATA <= x"38";
      when x"56A" => DATA <= x"A9";
      when x"56B" => DATA <= x"00";
      when x"56C" => DATA <= x"E5";
      when x"56D" => DATA <= x"6D";
      when x"56E" => DATA <= x"20";
      when x"56F" => DATA <= x"87";
      when x"570" => DATA <= x"D5";
      when x"571" => DATA <= x"A9";
      when x"572" => DATA <= x"0D";
      when x"573" => DATA <= x"D0";
      when x"574" => DATA <= x"18";
      when x"575" => DATA <= x"A5";
      when x"576" => DATA <= x"5A";
      when x"577" => DATA <= x"4A";
      when x"578" => DATA <= x"4A";
      when x"579" => DATA <= x"4A";
      when x"57A" => DATA <= x"4A";
      when x"57B" => DATA <= x"20";
      when x"57C" => DATA <= x"8B";
      when x"57D" => DATA <= x"D5";
      when x"57E" => DATA <= x"A5";
      when x"57F" => DATA <= x"5A";
      when x"580" => DATA <= x"29";
      when x"581" => DATA <= x"0F";
      when x"582" => DATA <= x"85";
      when x"583" => DATA <= x"5A";
      when x"584" => DATA <= x"4C";
      when x"585" => DATA <= x"4E";
      when x"586" => DATA <= x"D6";
      when x"587" => DATA <= x"C9";
      when x"588" => DATA <= x"0A";
      when x"589" => DATA <= x"B0";
      when x"58A" => DATA <= x"09";
      when x"58B" => DATA <= x"09";
      when x"58C" => DATA <= x"30";
      when x"58D" => DATA <= x"A4";
      when x"58E" => DATA <= x"6F";
      when x"58F" => DATA <= x"91";
      when x"590" => DATA <= x"52";
      when x"591" => DATA <= x"E6";
      when x"592" => DATA <= x"6F";
      when x"593" => DATA <= x"60";
      when x"594" => DATA <= x"A2";
      when x"595" => DATA <= x"FF";
      when x"596" => DATA <= x"E8";
      when x"597" => DATA <= x"E9";
      when x"598" => DATA <= x"0A";
      when x"599" => DATA <= x"B0";
      when x"59A" => DATA <= x"FB";
      when x"59B" => DATA <= x"69";
      when x"59C" => DATA <= x"0A";
      when x"59D" => DATA <= x"48";
      when x"59E" => DATA <= x"8A";
      when x"59F" => DATA <= x"20";
      when x"5A0" => DATA <= x"87";
      when x"5A1" => DATA <= x"D5";
      when x"5A2" => DATA <= x"68";
      when x"5A3" => DATA <= x"10";
      when x"5A4" => DATA <= x"E6";
      when x"5A5" => DATA <= x"A5";
      when x"5A6" => DATA <= x"03";
      when x"5A7" => DATA <= x"85";
      when x"5A8" => DATA <= x"54";
      when x"5A9" => DATA <= x"A5";
      when x"5AA" => DATA <= x"05";
      when x"5AB" => DATA <= x"85";
      when x"5AC" => DATA <= x"52";
      when x"5AD" => DATA <= x"A5";
      when x"5AE" => DATA <= x"06";
      when x"5AF" => DATA <= x"85";
      when x"5B0" => DATA <= x"53";
      when x"5B1" => DATA <= x"20";
      when x"5B2" => DATA <= x"A4";
      when x"5B3" => DATA <= x"DA";
      when x"5B4" => DATA <= x"85";
      when x"5B5" => DATA <= x"6C";
      when x"5B6" => DATA <= x"85";
      when x"5B7" => DATA <= x"6D";
      when x"5B8" => DATA <= x"20";
      when x"5B9" => DATA <= x"7B";
      when x"5BA" => DATA <= x"D6";
      when x"5BB" => DATA <= x"C9";
      when x"5BC" => DATA <= x"2E";
      when x"5BD" => DATA <= x"F0";
      when x"5BE" => DATA <= x"0E";
      when x"5BF" => DATA <= x"20";
      when x"5C0" => DATA <= x"C3";
      when x"5C1" => DATA <= x"D4";
      when x"5C2" => DATA <= x"90";
      when x"5C3" => DATA <= x"71";
      when x"5C4" => DATA <= x"85";
      when x"5C5" => DATA <= x"5E";
      when x"5C6" => DATA <= x"20";
      when x"5C7" => DATA <= x"7B";
      when x"5C8" => DATA <= x"D6";
      when x"5C9" => DATA <= x"C9";
      when x"5CA" => DATA <= x"2E";
      when x"5CB" => DATA <= x"D0";
      when x"5CC" => DATA <= x"09";
      when x"5CD" => DATA <= x"A5";
      when x"5CE" => DATA <= x"6C";
      when x"5CF" => DATA <= x"18";
      when x"5D0" => DATA <= x"D0";
      when x"5D1" => DATA <= x"3A";
      when x"5D2" => DATA <= x"E6";
      when x"5D3" => DATA <= x"6C";
      when x"5D4" => DATA <= x"D0";
      when x"5D5" => DATA <= x"F0";
      when x"5D6" => DATA <= x"C9";
      when x"5D7" => DATA <= x"45";
      when x"5D8" => DATA <= x"F0";
      when x"5D9" => DATA <= x"27";
      when x"5DA" => DATA <= x"20";
      when x"5DB" => DATA <= x"C3";
      when x"5DC" => DATA <= x"D4";
      when x"5DD" => DATA <= x"90";
      when x"5DE" => DATA <= x"2D";
      when x"5DF" => DATA <= x"85";
      when x"5E0" => DATA <= x"6E";
      when x"5E1" => DATA <= x"A5";
      when x"5E2" => DATA <= x"5A";
      when x"5E3" => DATA <= x"C9";
      when x"5E4" => DATA <= x"18";
      when x"5E5" => DATA <= x"90";
      when x"5E6" => DATA <= x"08";
      when x"5E7" => DATA <= x"A5";
      when x"5E8" => DATA <= x"6C";
      when x"5E9" => DATA <= x"D0";
      when x"5EA" => DATA <= x"DB";
      when x"5EB" => DATA <= x"E6";
      when x"5EC" => DATA <= x"6D";
      when x"5ED" => DATA <= x"B0";
      when x"5EE" => DATA <= x"D7";
      when x"5EF" => DATA <= x"A5";
      when x"5F0" => DATA <= x"6C";
      when x"5F1" => DATA <= x"F0";
      when x"5F2" => DATA <= x"02";
      when x"5F3" => DATA <= x"C6";
      when x"5F4" => DATA <= x"6D";
      when x"5F5" => DATA <= x"20";
      when x"5F6" => DATA <= x"4E";
      when x"5F7" => DATA <= x"D6";
      when x"5F8" => DATA <= x"18";
      when x"5F9" => DATA <= x"A5";
      when x"5FA" => DATA <= x"6E";
      when x"5FB" => DATA <= x"20";
      when x"5FC" => DATA <= x"36";
      when x"5FD" => DATA <= x"D6";
      when x"5FE" => DATA <= x"4C";
      when x"5FF" => DATA <= x"C6";
      when x"600" => DATA <= x"D5";
      when x"601" => DATA <= x"20";
      when x"602" => DATA <= x"7B";
      when x"603" => DATA <= x"D6";
      when x"604" => DATA <= x"20";
      when x"605" => DATA <= x"78";
      when x"606" => DATA <= x"D7";
      when x"607" => DATA <= x"18";
      when x"608" => DATA <= x"65";
      when x"609" => DATA <= x"6D";
      when x"60A" => DATA <= x"85";
      when x"60B" => DATA <= x"6D";
      when x"60C" => DATA <= x"A9";
      when x"60D" => DATA <= x"A8";
      when x"60E" => DATA <= x"85";
      when x"60F" => DATA <= x"59";
      when x"610" => DATA <= x"20";
      when x"611" => DATA <= x"86";
      when x"612" => DATA <= x"D6";
      when x"613" => DATA <= x"F0";
      when x"614" => DATA <= x"1C";
      when x"615" => DATA <= x"20";
      when x"616" => DATA <= x"C8";
      when x"617" => DATA <= x"D7";
      when x"618" => DATA <= x"A5";
      when x"619" => DATA <= x"6D";
      when x"61A" => DATA <= x"30";
      when x"61B" => DATA <= x"0B";
      when x"61C" => DATA <= x"F0";
      when x"61D" => DATA <= x"10";
      when x"61E" => DATA <= x"20";
      when x"61F" => DATA <= x"A0";
      when x"620" => DATA <= x"D6";
      when x"621" => DATA <= x"C6";
      when x"622" => DATA <= x"6D";
      when x"623" => DATA <= x"D0";
      when x"624" => DATA <= x"F9";
      when x"625" => DATA <= x"F0";
      when x"626" => DATA <= x"07";
      when x"627" => DATA <= x"20";
      when x"628" => DATA <= x"1B";
      when x"629" => DATA <= x"D7";
      when x"62A" => DATA <= x"E6";
      when x"62B" => DATA <= x"6D";
      when x"62C" => DATA <= x"D0";
      when x"62D" => DATA <= x"F9";
      when x"62E" => DATA <= x"20";
      when x"62F" => DATA <= x"9B";
      when x"630" => DATA <= x"DA";
      when x"631" => DATA <= x"38";
      when x"632" => DATA <= x"A4";
      when x"633" => DATA <= x"54";
      when x"634" => DATA <= x"88";
      when x"635" => DATA <= x"60";
      when x"636" => DATA <= x"A2";
      when x"637" => DATA <= x"05";
      when x"638" => DATA <= x"75";
      when x"639" => DATA <= x"59";
      when x"63A" => DATA <= x"95";
      when x"63B" => DATA <= x"59";
      when x"63C" => DATA <= x"A9";
      when x"63D" => DATA <= x"00";
      when x"63E" => DATA <= x"CA";
      when x"63F" => DATA <= x"D0";
      when x"640" => DATA <= x"F7";
      when x"641" => DATA <= x"60";
      when x"642" => DATA <= x"A2";
      when x"643" => DATA <= x"05";
      when x"644" => DATA <= x"B5";
      when x"645" => DATA <= x"59";
      when x"646" => DATA <= x"75";
      when x"647" => DATA <= x"61";
      when x"648" => DATA <= x"95";
      when x"649" => DATA <= x"59";
      when x"64A" => DATA <= x"CA";
      when x"64B" => DATA <= x"D0";
      when x"64C" => DATA <= x"F7";
      when x"64D" => DATA <= x"60";
      when x"64E" => DATA <= x"A2";
      when x"64F" => DATA <= x"05";
      when x"650" => DATA <= x"A9";
      when x"651" => DATA <= x"00";
      when x"652" => DATA <= x"85";
      when x"653" => DATA <= x"67";
      when x"654" => DATA <= x"A9";
      when x"655" => DATA <= x"00";
      when x"656" => DATA <= x"85";
      when x"657" => DATA <= x"68";
      when x"658" => DATA <= x"B5";
      when x"659" => DATA <= x"59";
      when x"65A" => DATA <= x"0A";
      when x"65B" => DATA <= x"26";
      when x"65C" => DATA <= x"68";
      when x"65D" => DATA <= x"0A";
      when x"65E" => DATA <= x"26";
      when x"65F" => DATA <= x"68";
      when x"660" => DATA <= x"18";
      when x"661" => DATA <= x"75";
      when x"662" => DATA <= x"59";
      when x"663" => DATA <= x"90";
      when x"664" => DATA <= x"02";
      when x"665" => DATA <= x"E6";
      when x"666" => DATA <= x"68";
      when x"667" => DATA <= x"0A";
      when x"668" => DATA <= x"26";
      when x"669" => DATA <= x"68";
      when x"66A" => DATA <= x"18";
      when x"66B" => DATA <= x"65";
      when x"66C" => DATA <= x"67";
      when x"66D" => DATA <= x"90";
      when x"66E" => DATA <= x"02";
      when x"66F" => DATA <= x"E6";
      when x"670" => DATA <= x"68";
      when x"671" => DATA <= x"95";
      when x"672" => DATA <= x"59";
      when x"673" => DATA <= x"A5";
      when x"674" => DATA <= x"68";
      when x"675" => DATA <= x"85";
      when x"676" => DATA <= x"67";
      when x"677" => DATA <= x"CA";
      when x"678" => DATA <= x"D0";
      when x"679" => DATA <= x"DA";
      when x"67A" => DATA <= x"60";
      when x"67B" => DATA <= x"84";
      when x"67C" => DATA <= x"55";
      when x"67D" => DATA <= x"A4";
      when x"67E" => DATA <= x"54";
      when x"67F" => DATA <= x"B1";
      when x"680" => DATA <= x"52";
      when x"681" => DATA <= x"A4";
      when x"682" => DATA <= x"55";
      when x"683" => DATA <= x"E6";
      when x"684" => DATA <= x"54";
      when x"685" => DATA <= x"60";
      when x"686" => DATA <= x"A5";
      when x"687" => DATA <= x"5A";
      when x"688" => DATA <= x"05";
      when x"689" => DATA <= x"5B";
      when x"68A" => DATA <= x"05";
      when x"68B" => DATA <= x"5C";
      when x"68C" => DATA <= x"05";
      when x"68D" => DATA <= x"5D";
      when x"68E" => DATA <= x"05";
      when x"68F" => DATA <= x"5E";
      when x"690" => DATA <= x"F0";
      when x"691" => DATA <= x"07";
      when x"692" => DATA <= x"A5";
      when x"693" => DATA <= x"57";
      when x"694" => DATA <= x"D0";
      when x"695" => DATA <= x"09";
      when x"696" => DATA <= x"A9";
      when x"697" => DATA <= x"01";
      when x"698" => DATA <= x"60";
      when x"699" => DATA <= x"85";
      when x"69A" => DATA <= x"57";
      when x"69B" => DATA <= x"85";
      when x"69C" => DATA <= x"59";
      when x"69D" => DATA <= x"85";
      when x"69E" => DATA <= x"58";
      when x"69F" => DATA <= x"60";
      when x"6A0" => DATA <= x"18";
      when x"6A1" => DATA <= x"A5";
      when x"6A2" => DATA <= x"59";
      when x"6A3" => DATA <= x"69";
      when x"6A4" => DATA <= x"03";
      when x"6A5" => DATA <= x"85";
      when x"6A6" => DATA <= x"59";
      when x"6A7" => DATA <= x"90";
      when x"6A8" => DATA <= x"02";
      when x"6A9" => DATA <= x"E6";
      when x"6AA" => DATA <= x"58";
      when x"6AB" => DATA <= x"20";
      when x"6AC" => DATA <= x"C3";
      when x"6AD" => DATA <= x"D6";
      when x"6AE" => DATA <= x"20";
      when x"6AF" => DATA <= x"FB";
      when x"6B0" => DATA <= x"D6";
      when x"6B1" => DATA <= x"20";
      when x"6B2" => DATA <= x"FB";
      when x"6B3" => DATA <= x"D6";
      when x"6B4" => DATA <= x"20";
      when x"6B5" => DATA <= x"42";
      when x"6B6" => DATA <= x"D6";
      when x"6B7" => DATA <= x"90";
      when x"6B8" => DATA <= x"09";
      when x"6B9" => DATA <= x"20";
      when x"6BA" => DATA <= x"D8";
      when x"6BB" => DATA <= x"D6";
      when x"6BC" => DATA <= x"E6";
      when x"6BD" => DATA <= x"59";
      when x"6BE" => DATA <= x"D0";
      when x"6BF" => DATA <= x"02";
      when x"6C0" => DATA <= x"E6";
      when x"6C1" => DATA <= x"58";
      when x"6C2" => DATA <= x"60";
      when x"6C3" => DATA <= x"A2";
      when x"6C4" => DATA <= x"08";
      when x"6C5" => DATA <= x"B5";
      when x"6C6" => DATA <= x"56";
      when x"6C7" => DATA <= x"95";
      when x"6C8" => DATA <= x"5E";
      when x"6C9" => DATA <= x"CA";
      when x"6CA" => DATA <= x"D0";
      when x"6CB" => DATA <= x"F9";
      when x"6CC" => DATA <= x"60";
      when x"6CD" => DATA <= x"06";
      when x"6CE" => DATA <= x"5E";
      when x"6CF" => DATA <= x"26";
      when x"6D0" => DATA <= x"5D";
      when x"6D1" => DATA <= x"26";
      when x"6D2" => DATA <= x"5C";
      when x"6D3" => DATA <= x"26";
      when x"6D4" => DATA <= x"5B";
      when x"6D5" => DATA <= x"26";
      when x"6D6" => DATA <= x"5A";
      when x"6D7" => DATA <= x"60";
      when x"6D8" => DATA <= x"66";
      when x"6D9" => DATA <= x"5A";
      when x"6DA" => DATA <= x"66";
      when x"6DB" => DATA <= x"5B";
      when x"6DC" => DATA <= x"66";
      when x"6DD" => DATA <= x"5C";
      when x"6DE" => DATA <= x"66";
      when x"6DF" => DATA <= x"5D";
      when x"6E0" => DATA <= x"66";
      when x"6E1" => DATA <= x"5E";
      when x"6E2" => DATA <= x"60";
      when x"6E3" => DATA <= x"A5";
      when x"6E4" => DATA <= x"5D";
      when x"6E5" => DATA <= x"85";
      when x"6E6" => DATA <= x"5E";
      when x"6E7" => DATA <= x"A5";
      when x"6E8" => DATA <= x"5C";
      when x"6E9" => DATA <= x"85";
      when x"6EA" => DATA <= x"5D";
      when x"6EB" => DATA <= x"A5";
      when x"6EC" => DATA <= x"5B";
      when x"6ED" => DATA <= x"85";
      when x"6EE" => DATA <= x"5C";
      when x"6EF" => DATA <= x"A5";
      when x"6F0" => DATA <= x"5A";
      when x"6F1" => DATA <= x"85";
      when x"6F2" => DATA <= x"5B";
      when x"6F3" => DATA <= x"A9";
      when x"6F4" => DATA <= x"00";
      when x"6F5" => DATA <= x"85";
      when x"6F6" => DATA <= x"5A";
      when x"6F7" => DATA <= x"60";
      when x"6F8" => DATA <= x"20";
      when x"6F9" => DATA <= x"C3";
      when x"6FA" => DATA <= x"D6";
      when x"6FB" => DATA <= x"46";
      when x"6FC" => DATA <= x"62";
      when x"6FD" => DATA <= x"66";
      when x"6FE" => DATA <= x"63";
      when x"6FF" => DATA <= x"66";
      when x"700" => DATA <= x"64";
      when x"701" => DATA <= x"66";
      when x"702" => DATA <= x"65";
      when x"703" => DATA <= x"66";
      when x"704" => DATA <= x"66";
      when x"705" => DATA <= x"60";
      when x"706" => DATA <= x"A5";
      when x"707" => DATA <= x"65";
      when x"708" => DATA <= x"85";
      when x"709" => DATA <= x"66";
      when x"70A" => DATA <= x"A5";
      when x"70B" => DATA <= x"64";
      when x"70C" => DATA <= x"85";
      when x"70D" => DATA <= x"65";
      when x"70E" => DATA <= x"A5";
      when x"70F" => DATA <= x"63";
      when x"710" => DATA <= x"85";
      when x"711" => DATA <= x"64";
      when x"712" => DATA <= x"A5";
      when x"713" => DATA <= x"62";
      when x"714" => DATA <= x"85";
      when x"715" => DATA <= x"63";
      when x"716" => DATA <= x"A9";
      when x"717" => DATA <= x"00";
      when x"718" => DATA <= x"85";
      when x"719" => DATA <= x"62";
      when x"71A" => DATA <= x"60";
      when x"71B" => DATA <= x"38";
      when x"71C" => DATA <= x"A5";
      when x"71D" => DATA <= x"59";
      when x"71E" => DATA <= x"E9";
      when x"71F" => DATA <= x"04";
      when x"720" => DATA <= x"85";
      when x"721" => DATA <= x"59";
      when x"722" => DATA <= x"B0";
      when x"723" => DATA <= x"02";
      when x"724" => DATA <= x"C6";
      when x"725" => DATA <= x"58";
      when x"726" => DATA <= x"20";
      when x"727" => DATA <= x"F8";
      when x"728" => DATA <= x"D6";
      when x"729" => DATA <= x"20";
      when x"72A" => DATA <= x"B4";
      when x"72B" => DATA <= x"D6";
      when x"72C" => DATA <= x"20";
      when x"72D" => DATA <= x"F8";
      when x"72E" => DATA <= x"D6";
      when x"72F" => DATA <= x"20";
      when x"730" => DATA <= x"FB";
      when x"731" => DATA <= x"D6";
      when x"732" => DATA <= x"20";
      when x"733" => DATA <= x"FB";
      when x"734" => DATA <= x"D6";
      when x"735" => DATA <= x"20";
      when x"736" => DATA <= x"FB";
      when x"737" => DATA <= x"D6";
      when x"738" => DATA <= x"20";
      when x"739" => DATA <= x"B4";
      when x"73A" => DATA <= x"D6";
      when x"73B" => DATA <= x"A9";
      when x"73C" => DATA <= x"00";
      when x"73D" => DATA <= x"85";
      when x"73E" => DATA <= x"62";
      when x"73F" => DATA <= x"A5";
      when x"740" => DATA <= x"5A";
      when x"741" => DATA <= x"85";
      when x"742" => DATA <= x"63";
      when x"743" => DATA <= x"A5";
      when x"744" => DATA <= x"5B";
      when x"745" => DATA <= x"85";
      when x"746" => DATA <= x"64";
      when x"747" => DATA <= x"A5";
      when x"748" => DATA <= x"5C";
      when x"749" => DATA <= x"85";
      when x"74A" => DATA <= x"65";
      when x"74B" => DATA <= x"A5";
      when x"74C" => DATA <= x"5D";
      when x"74D" => DATA <= x"85";
      when x"74E" => DATA <= x"66";
      when x"74F" => DATA <= x"A5";
      when x"750" => DATA <= x"5E";
      when x"751" => DATA <= x"2A";
      when x"752" => DATA <= x"20";
      when x"753" => DATA <= x"B4";
      when x"754" => DATA <= x"D6";
      when x"755" => DATA <= x"A9";
      when x"756" => DATA <= x"00";
      when x"757" => DATA <= x"85";
      when x"758" => DATA <= x"62";
      when x"759" => DATA <= x"85";
      when x"75A" => DATA <= x"63";
      when x"75B" => DATA <= x"A5";
      when x"75C" => DATA <= x"5A";
      when x"75D" => DATA <= x"85";
      when x"75E" => DATA <= x"64";
      when x"75F" => DATA <= x"A5";
      when x"760" => DATA <= x"5B";
      when x"761" => DATA <= x"85";
      when x"762" => DATA <= x"65";
      when x"763" => DATA <= x"A5";
      when x"764" => DATA <= x"5C";
      when x"765" => DATA <= x"85";
      when x"766" => DATA <= x"66";
      when x"767" => DATA <= x"A5";
      when x"768" => DATA <= x"5D";
      when x"769" => DATA <= x"2A";
      when x"76A" => DATA <= x"20";
      when x"76B" => DATA <= x"B4";
      when x"76C" => DATA <= x"D6";
      when x"76D" => DATA <= x"A5";
      when x"76E" => DATA <= x"5B";
      when x"76F" => DATA <= x"2A";
      when x"770" => DATA <= x"A5";
      when x"771" => DATA <= x"5A";
      when x"772" => DATA <= x"20";
      when x"773" => DATA <= x"36";
      when x"774" => DATA <= x"D6";
      when x"775" => DATA <= x"4C";
      when x"776" => DATA <= x"B7";
      when x"777" => DATA <= x"D6";
      when x"778" => DATA <= x"A0";
      when x"779" => DATA <= x"FF";
      when x"77A" => DATA <= x"C9";
      when x"77B" => DATA <= x"2B";
      when x"77C" => DATA <= x"F0";
      when x"77D" => DATA <= x"05";
      when x"77E" => DATA <= x"C9";
      when x"77F" => DATA <= x"2D";
      when x"780" => DATA <= x"D0";
      when x"781" => DATA <= x"04";
      when x"782" => DATA <= x"C8";
      when x"783" => DATA <= x"20";
      when x"784" => DATA <= x"7B";
      when x"785" => DATA <= x"D6";
      when x"786" => DATA <= x"20";
      when x"787" => DATA <= x"C3";
      when x"788" => DATA <= x"D4";
      when x"789" => DATA <= x"90";
      when x"78A" => DATA <= x"24";
      when x"78B" => DATA <= x"AA";
      when x"78C" => DATA <= x"20";
      when x"78D" => DATA <= x"7B";
      when x"78E" => DATA <= x"D6";
      when x"78F" => DATA <= x"20";
      when x"790" => DATA <= x"C3";
      when x"791" => DATA <= x"D4";
      when x"792" => DATA <= x"90";
      when x"793" => DATA <= x"10";
      when x"794" => DATA <= x"85";
      when x"795" => DATA <= x"6E";
      when x"796" => DATA <= x"20";
      when x"797" => DATA <= x"7B";
      when x"798" => DATA <= x"D6";
      when x"799" => DATA <= x"8A";
      when x"79A" => DATA <= x"85";
      when x"79B" => DATA <= x"67";
      when x"79C" => DATA <= x"0A";
      when x"79D" => DATA <= x"0A";
      when x"79E" => DATA <= x"65";
      when x"79F" => DATA <= x"67";
      when x"7A0" => DATA <= x"0A";
      when x"7A1" => DATA <= x"65";
      when x"7A2" => DATA <= x"6E";
      when x"7A3" => DATA <= x"AA";
      when x"7A4" => DATA <= x"98";
      when x"7A5" => DATA <= x"D0";
      when x"7A6" => DATA <= x"06";
      when x"7A7" => DATA <= x"86";
      when x"7A8" => DATA <= x"6E";
      when x"7A9" => DATA <= x"38";
      when x"7AA" => DATA <= x"E5";
      when x"7AB" => DATA <= x"6E";
      when x"7AC" => DATA <= x"60";
      when x"7AD" => DATA <= x"8A";
      when x"7AE" => DATA <= x"60";
      when x"7AF" => DATA <= x"A9";
      when x"7B0" => DATA <= x"00";
      when x"7B1" => DATA <= x"60";
      when x"7B2" => DATA <= x"48";
      when x"7B3" => DATA <= x"20";
      when x"7B4" => DATA <= x"A4";
      when x"7B5" => DATA <= x"DA";
      when x"7B6" => DATA <= x"68";
      when x"7B7" => DATA <= x"F0";
      when x"7B8" => DATA <= x"F8";
      when x"7B9" => DATA <= x"10";
      when x"7BA" => DATA <= x"07";
      when x"7BB" => DATA <= x"85";
      when x"7BC" => DATA <= x"57";
      when x"7BD" => DATA <= x"A9";
      when x"7BE" => DATA <= x"00";
      when x"7BF" => DATA <= x"38";
      when x"7C0" => DATA <= x"E5";
      when x"7C1" => DATA <= x"57";
      when x"7C2" => DATA <= x"85";
      when x"7C3" => DATA <= x"5A";
      when x"7C4" => DATA <= x"A9";
      when x"7C5" => DATA <= x"88";
      when x"7C6" => DATA <= x"85";
      when x"7C7" => DATA <= x"59";
      when x"7C8" => DATA <= x"20";
      when x"7C9" => DATA <= x"86";
      when x"7CA" => DATA <= x"D6";
      when x"7CB" => DATA <= x"F0";
      when x"7CC" => DATA <= x"E4";
      when x"7CD" => DATA <= x"A5";
      when x"7CE" => DATA <= x"5A";
      when x"7CF" => DATA <= x"D0";
      when x"7D0" => DATA <= x"21";
      when x"7D1" => DATA <= x"A5";
      when x"7D2" => DATA <= x"5B";
      when x"7D3" => DATA <= x"85";
      when x"7D4" => DATA <= x"5A";
      when x"7D5" => DATA <= x"A5";
      when x"7D6" => DATA <= x"5C";
      when x"7D7" => DATA <= x"85";
      when x"7D8" => DATA <= x"5B";
      when x"7D9" => DATA <= x"A5";
      when x"7DA" => DATA <= x"5D";
      when x"7DB" => DATA <= x"85";
      when x"7DC" => DATA <= x"5C";
      when x"7DD" => DATA <= x"A5";
      when x"7DE" => DATA <= x"5E";
      when x"7DF" => DATA <= x"85";
      when x"7E0" => DATA <= x"5D";
      when x"7E1" => DATA <= x"A9";
      when x"7E2" => DATA <= x"00";
      when x"7E3" => DATA <= x"85";
      when x"7E4" => DATA <= x"5E";
      when x"7E5" => DATA <= x"38";
      when x"7E6" => DATA <= x"A5";
      when x"7E7" => DATA <= x"59";
      when x"7E8" => DATA <= x"E9";
      when x"7E9" => DATA <= x"08";
      when x"7EA" => DATA <= x"85";
      when x"7EB" => DATA <= x"59";
      when x"7EC" => DATA <= x"B0";
      when x"7ED" => DATA <= x"DF";
      when x"7EE" => DATA <= x"C6";
      when x"7EF" => DATA <= x"58";
      when x"7F0" => DATA <= x"90";
      when x"7F1" => DATA <= x"DB";
      when x"7F2" => DATA <= x"A5";
      when x"7F3" => DATA <= x"5A";
      when x"7F4" => DATA <= x"30";
      when x"7F5" => DATA <= x"BB";
      when x"7F6" => DATA <= x"20";
      when x"7F7" => DATA <= x"CD";
      when x"7F8" => DATA <= x"D6";
      when x"7F9" => DATA <= x"A5";
      when x"7FA" => DATA <= x"59";
      when x"7FB" => DATA <= x"D0";
      when x"7FC" => DATA <= x"02";
      when x"7FD" => DATA <= x"C6";
      when x"7FE" => DATA <= x"58";
      when x"7FF" => DATA <= x"C6";
      when x"800" => DATA <= x"59";
      when x"801" => DATA <= x"4C";
      when x"802" => DATA <= x"F2";
      when x"803" => DATA <= x"D7";
      when x"804" => DATA <= x"A0";
      when x"805" => DATA <= x"04";
      when x"806" => DATA <= x"A9";
      when x"807" => DATA <= x"00";
      when x"808" => DATA <= x"85";
      when x"809" => DATA <= x"66";
      when x"80A" => DATA <= x"85";
      when x"80B" => DATA <= x"60";
      when x"80C" => DATA <= x"85";
      when x"80D" => DATA <= x"5F";
      when x"80E" => DATA <= x"B1";
      when x"80F" => DATA <= x"6F";
      when x"810" => DATA <= x"99";
      when x"811" => DATA <= x"61";
      when x"812" => DATA <= x"00";
      when x"813" => DATA <= x"05";
      when x"814" => DATA <= x"5F";
      when x"815" => DATA <= x"85";
      when x"816" => DATA <= x"5F";
      when x"817" => DATA <= x"88";
      when x"818" => DATA <= x"10";
      when x"819" => DATA <= x"F4";
      when x"81A" => DATA <= x"AA";
      when x"81B" => DATA <= x"F0";
      when x"81C" => DATA <= x"09";
      when x"81D" => DATA <= x"A5";
      when x"81E" => DATA <= x"62";
      when x"81F" => DATA <= x"85";
      when x"820" => DATA <= x"5F";
      when x"821" => DATA <= x"09";
      when x"822" => DATA <= x"80";
      when x"823" => DATA <= x"85";
      when x"824" => DATA <= x"62";
      when x"825" => DATA <= x"8A";
      when x"826" => DATA <= x"60";
      when x"827" => DATA <= x"20";
      when x"828" => DATA <= x"A2";
      when x"829" => DATA <= x"DB";
      when x"82A" => DATA <= x"D0";
      when x"82B" => DATA <= x"11";
      when x"82C" => DATA <= x"20";
      when x"82D" => DATA <= x"A6";
      when x"82E" => DATA <= x"DB";
      when x"82F" => DATA <= x"D0";
      when x"830" => DATA <= x"0C";
      when x"831" => DATA <= x"20";
      when x"832" => DATA <= x"AA";
      when x"833" => DATA <= x"DB";
      when x"834" => DATA <= x"D0";
      when x"835" => DATA <= x"07";
      when x"836" => DATA <= x"A6";
      when x"837" => DATA <= x"04";
      when x"838" => DATA <= x"A0";
      when x"839" => DATA <= x"6F";
      when x"83A" => DATA <= x"20";
      when x"83B" => DATA <= x"CD";
      when x"83C" => DATA <= x"C3";
      when x"83D" => DATA <= x"A0";
      when x"83E" => DATA <= x"00";
      when x"83F" => DATA <= x"A5";
      when x"840" => DATA <= x"59";
      when x"841" => DATA <= x"91";
      when x"842" => DATA <= x"6F";
      when x"843" => DATA <= x"C8";
      when x"844" => DATA <= x"A5";
      when x"845" => DATA <= x"57";
      when x"846" => DATA <= x"29";
      when x"847" => DATA <= x"80";
      when x"848" => DATA <= x"85";
      when x"849" => DATA <= x"57";
      when x"84A" => DATA <= x"A5";
      when x"84B" => DATA <= x"5A";
      when x"84C" => DATA <= x"29";
      when x"84D" => DATA <= x"7F";
      when x"84E" => DATA <= x"05";
      when x"84F" => DATA <= x"57";
      when x"850" => DATA <= x"91";
      when x"851" => DATA <= x"6F";
      when x"852" => DATA <= x"C8";
      when x"853" => DATA <= x"B9";
      when x"854" => DATA <= x"59";
      when x"855" => DATA <= x"00";
      when x"856" => DATA <= x"91";
      when x"857" => DATA <= x"6F";
      when x"858" => DATA <= x"C0";
      when x"859" => DATA <= x"04";
      when x"85A" => DATA <= x"D0";
      when x"85B" => DATA <= x"F6";
      when x"85C" => DATA <= x"60";
      when x"85D" => DATA <= x"A0";
      when x"85E" => DATA <= x"52";
      when x"85F" => DATA <= x"84";
      when x"860" => DATA <= x"6F";
      when x"861" => DATA <= x"A9";
      when x"862" => DATA <= x"00";
      when x"863" => DATA <= x"85";
      when x"864" => DATA <= x"70";
      when x"865" => DATA <= x"20";
      when x"866" => DATA <= x"3D";
      when x"867" => DATA <= x"D8";
      when x"868" => DATA <= x"20";
      when x"869" => DATA <= x"D9";
      when x"86A" => DATA <= x"C4";
      when x"86B" => DATA <= x"A5";
      when x"86C" => DATA <= x"56";
      when x"86D" => DATA <= x"95";
      when x"86E" => DATA <= x"73";
      when x"86F" => DATA <= x"60";
      when x"870" => DATA <= x"A6";
      when x"871" => DATA <= x"04";
      when x"872" => DATA <= x"20";
      when x"873" => DATA <= x"CB";
      when x"874" => DATA <= x"C3";
      when x"875" => DATA <= x"B5";
      when x"876" => DATA <= x"74";
      when x"877" => DATA <= x"85";
      when x"878" => DATA <= x"56";
      when x"879" => DATA <= x"84";
      when x"87A" => DATA <= x"6F";
      when x"87B" => DATA <= x"A9";
      when x"87C" => DATA <= x"00";
      when x"87D" => DATA <= x"85";
      when x"87E" => DATA <= x"70";
      when x"87F" => DATA <= x"60";
      when x"880" => DATA <= x"A5";
      when x"881" => DATA <= x"5E";
      when x"882" => DATA <= x"C9";
      when x"883" => DATA <= x"80";
      when x"884" => DATA <= x"90";
      when x"885" => DATA <= x"07";
      when x"886" => DATA <= x"F0";
      when x"887" => DATA <= x"0A";
      when x"888" => DATA <= x"A9";
      when x"889" => DATA <= x"FF";
      when x"88A" => DATA <= x"20";
      when x"88B" => DATA <= x"72";
      when x"88C" => DATA <= x"D7";
      when x"88D" => DATA <= x"A9";
      when x"88E" => DATA <= x"00";
      when x"88F" => DATA <= x"85";
      when x"890" => DATA <= x"5E";
      when x"891" => DATA <= x"60";
      when x"892" => DATA <= x"A5";
      when x"893" => DATA <= x"5D";
      when x"894" => DATA <= x"09";
      when x"895" => DATA <= x"01";
      when x"896" => DATA <= x"85";
      when x"897" => DATA <= x"5D";
      when x"898" => DATA <= x"D0";
      when x"899" => DATA <= x"F3";
      when x"89A" => DATA <= x"20";
      when x"89B" => DATA <= x"C7";
      when x"89C" => DATA <= x"D8";
      when x"89D" => DATA <= x"F0";
      when x"89E" => DATA <= x"06";
      when x"89F" => DATA <= x"A5";
      when x"8A0" => DATA <= x"59";
      when x"8A1" => DATA <= x"C9";
      when x"8A2" => DATA <= x"A0";
      when x"8A3" => DATA <= x"B0";
      when x"8A4" => DATA <= x"14";
      when x"8A5" => DATA <= x"46";
      when x"8A6" => DATA <= x"5A";
      when x"8A7" => DATA <= x"66";
      when x"8A8" => DATA <= x"5B";
      when x"8A9" => DATA <= x"66";
      when x"8AA" => DATA <= x"5C";
      when x"8AB" => DATA <= x"66";
      when x"8AC" => DATA <= x"5D";
      when x"8AD" => DATA <= x"66";
      when x"8AE" => DATA <= x"62";
      when x"8AF" => DATA <= x"66";
      when x"8B0" => DATA <= x"63";
      when x"8B1" => DATA <= x"66";
      when x"8B2" => DATA <= x"64";
      when x"8B3" => DATA <= x"66";
      when x"8B4" => DATA <= x"65";
      when x"8B5" => DATA <= x"E6";
      when x"8B6" => DATA <= x"59";
      when x"8B7" => DATA <= x"D0";
      when x"8B8" => DATA <= x"E6";
      when x"8B9" => DATA <= x"F0";
      when x"8BA" => DATA <= x"16";
      when x"8BB" => DATA <= x"A9";
      when x"8BC" => DATA <= x"7F";
      when x"8BD" => DATA <= x"85";
      when x"8BE" => DATA <= x"5A";
      when x"8BF" => DATA <= x"A9";
      when x"8C0" => DATA <= x"FF";
      when x"8C1" => DATA <= x"85";
      when x"8C2" => DATA <= x"5B";
      when x"8C3" => DATA <= x"85";
      when x"8C4" => DATA <= x"5C";
      when x"8C5" => DATA <= x"85";
      when x"8C6" => DATA <= x"5D";
      when x"8C7" => DATA <= x"A2";
      when x"8C8" => DATA <= x"08";
      when x"8C9" => DATA <= x"A9";
      when x"8CA" => DATA <= x"00";
      when x"8CB" => DATA <= x"95";
      when x"8CC" => DATA <= x"5F";
      when x"8CD" => DATA <= x"CA";
      when x"8CE" => DATA <= x"D0";
      when x"8CF" => DATA <= x"FB";
      when x"8D0" => DATA <= x"60";
      when x"8D1" => DATA <= x"A5";
      when x"8D2" => DATA <= x"57";
      when x"8D3" => DATA <= x"10";
      when x"8D4" => DATA <= x"0C";
      when x"8D5" => DATA <= x"38";
      when x"8D6" => DATA <= x"A2";
      when x"8D7" => DATA <= x"04";
      when x"8D8" => DATA <= x"A9";
      when x"8D9" => DATA <= x"00";
      when x"8DA" => DATA <= x"F5";
      when x"8DB" => DATA <= x"59";
      when x"8DC" => DATA <= x"95";
      when x"8DD" => DATA <= x"59";
      when x"8DE" => DATA <= x"CA";
      when x"8DF" => DATA <= x"D0";
      when x"8E0" => DATA <= x"F7";
      when x"8E1" => DATA <= x"60";
      when x"8E2" => DATA <= x"A5";
      when x"8E3" => DATA <= x"62";
      when x"8E4" => DATA <= x"10";
      when x"8E5" => DATA <= x"23";
      when x"8E6" => DATA <= x"A2";
      when x"8E7" => DATA <= x"04";
      when x"8E8" => DATA <= x"A9";
      when x"8E9" => DATA <= x"00";
      when x"8EA" => DATA <= x"F5";
      when x"8EB" => DATA <= x"61";
      when x"8EC" => DATA <= x"95";
      when x"8ED" => DATA <= x"61";
      when x"8EE" => DATA <= x"CA";
      when x"8EF" => DATA <= x"D0";
      when x"8F0" => DATA <= x"F7";
      when x"8F1" => DATA <= x"A5";
      when x"8F2" => DATA <= x"57";
      when x"8F3" => DATA <= x"49";
      when x"8F4" => DATA <= x"80";
      when x"8F5" => DATA <= x"85";
      when x"8F6" => DATA <= x"57";
      when x"8F7" => DATA <= x"10";
      when x"8F8" => DATA <= x"11";
      when x"8F9" => DATA <= x"E6";
      when x"8FA" => DATA <= x"5D";
      when x"8FB" => DATA <= x"D0";
      when x"8FC" => DATA <= x"0C";
      when x"8FD" => DATA <= x"E6";
      when x"8FE" => DATA <= x"5C";
      when x"8FF" => DATA <= x"D0";
      when x"900" => DATA <= x"08";
      when x"901" => DATA <= x"E6";
      when x"902" => DATA <= x"5B";
      when x"903" => DATA <= x"D0";
      when x"904" => DATA <= x"04";
      when x"905" => DATA <= x"E6";
      when x"906" => DATA <= x"5A";
      when x"907" => DATA <= x"F0";
      when x"908" => DATA <= x"B2";
      when x"909" => DATA <= x"60";
      when x"90A" => DATA <= x"20";
      when x"90B" => DATA <= x"D5";
      when x"90C" => DATA <= x"D8";
      when x"90D" => DATA <= x"20";
      when x"90E" => DATA <= x"F9";
      when x"90F" => DATA <= x"D8";
      when x"910" => DATA <= x"4C";
      when x"911" => DATA <= x"D5";
      when x"912" => DATA <= x"D8";
      when x"913" => DATA <= x"A2";
      when x"914" => DATA <= x"05";
      when x"915" => DATA <= x"B5";
      when x"916" => DATA <= x"61";
      when x"917" => DATA <= x"95";
      when x"918" => DATA <= x"59";
      when x"919" => DATA <= x"CA";
      when x"91A" => DATA <= x"D0";
      when x"91B" => DATA <= x"F9";
      when x"91C" => DATA <= x"A9";
      when x"91D" => DATA <= x"80";
      when x"91E" => DATA <= x"85";
      when x"91F" => DATA <= x"59";
      when x"920" => DATA <= x"4C";
      when x"921" => DATA <= x"C8";
      when x"922" => DATA <= x"D7";
      when x"923" => DATA <= x"20";
      when x"924" => DATA <= x"04";
      when x"925" => DATA <= x"D8";
      when x"926" => DATA <= x"20";
      when x"927" => DATA <= x"3D";
      when x"928" => DATA <= x"D8";
      when x"929" => DATA <= x"A2";
      when x"92A" => DATA <= x"08";
      when x"92B" => DATA <= x"B5";
      when x"92C" => DATA <= x"5E";
      when x"92D" => DATA <= x"95";
      when x"92E" => DATA <= x"56";
      when x"92F" => DATA <= x"CA";
      when x"930" => DATA <= x"D0";
      when x"931" => DATA <= x"F9";
      when x"932" => DATA <= x"60";
      when x"933" => DATA <= x"20";
      when x"934" => DATA <= x"39";
      when x"935" => DATA <= x"D9";
      when x"936" => DATA <= x"4C";
      when x"937" => DATA <= x"BF";
      when x"938" => DATA <= x"D1";
      when x"939" => DATA <= x"20";
      when x"93A" => DATA <= x"BF";
      when x"93B" => DATA <= x"D1";
      when x"93C" => DATA <= x"20";
      when x"93D" => DATA <= x"04";
      when x"93E" => DATA <= x"D8";
      when x"93F" => DATA <= x"F0";
      when x"940" => DATA <= x"F1";
      when x"941" => DATA <= x"20";
      when x"942" => DATA <= x"86";
      when x"943" => DATA <= x"D6";
      when x"944" => DATA <= x"F0";
      when x"945" => DATA <= x"E3";
      when x"946" => DATA <= x"A5";
      when x"947" => DATA <= x"59";
      when x"948" => DATA <= x"C5";
      when x"949" => DATA <= x"61";
      when x"94A" => DATA <= x"F0";
      when x"94B" => DATA <= x"26";
      when x"94C" => DATA <= x"90";
      when x"94D" => DATA <= x"0F";
      when x"94E" => DATA <= x"E5";
      when x"94F" => DATA <= x"61";
      when x"950" => DATA <= x"C9";
      when x"951" => DATA <= x"21";
      when x"952" => DATA <= x"B0";
      when x"953" => DATA <= x"DE";
      when x"954" => DATA <= x"AA";
      when x"955" => DATA <= x"20";
      when x"956" => DATA <= x"FB";
      when x"957" => DATA <= x"D6";
      when x"958" => DATA <= x"CA";
      when x"959" => DATA <= x"D0";
      when x"95A" => DATA <= x"FA";
      when x"95B" => DATA <= x"F0";
      when x"95C" => DATA <= x"15";
      when x"95D" => DATA <= x"38";
      when x"95E" => DATA <= x"A5";
      when x"95F" => DATA <= x"61";
      when x"960" => DATA <= x"E5";
      when x"961" => DATA <= x"59";
      when x"962" => DATA <= x"C9";
      when x"963" => DATA <= x"21";
      when x"964" => DATA <= x"B0";
      when x"965" => DATA <= x"C3";
      when x"966" => DATA <= x"AA";
      when x"967" => DATA <= x"18";
      when x"968" => DATA <= x"20";
      when x"969" => DATA <= x"D8";
      when x"96A" => DATA <= x"D6";
      when x"96B" => DATA <= x"CA";
      when x"96C" => DATA <= x"D0";
      when x"96D" => DATA <= x"F9";
      when x"96E" => DATA <= x"A5";
      when x"96F" => DATA <= x"61";
      when x"970" => DATA <= x"85";
      when x"971" => DATA <= x"59";
      when x"972" => DATA <= x"A5";
      when x"973" => DATA <= x"57";
      when x"974" => DATA <= x"45";
      when x"975" => DATA <= x"5F";
      when x"976" => DATA <= x"10";
      when x"977" => DATA <= x"49";
      when x"978" => DATA <= x"A5";
      when x"979" => DATA <= x"5A";
      when x"97A" => DATA <= x"C5";
      when x"97B" => DATA <= x"62";
      when x"97C" => DATA <= x"D0";
      when x"97D" => DATA <= x"1B";
      when x"97E" => DATA <= x"A5";
      when x"97F" => DATA <= x"5B";
      when x"980" => DATA <= x"C5";
      when x"981" => DATA <= x"63";
      when x"982" => DATA <= x"D0";
      when x"983" => DATA <= x"15";
      when x"984" => DATA <= x"A5";
      when x"985" => DATA <= x"5C";
      when x"986" => DATA <= x"C5";
      when x"987" => DATA <= x"64";
      when x"988" => DATA <= x"D0";
      when x"989" => DATA <= x"0F";
      when x"98A" => DATA <= x"A5";
      when x"98B" => DATA <= x"5D";
      when x"98C" => DATA <= x"C5";
      when x"98D" => DATA <= x"65";
      when x"98E" => DATA <= x"D0";
      when x"98F" => DATA <= x"09";
      when x"990" => DATA <= x"A5";
      when x"991" => DATA <= x"5E";
      when x"992" => DATA <= x"C5";
      when x"993" => DATA <= x"66";
      when x"994" => DATA <= x"D0";
      when x"995" => DATA <= x"03";
      when x"996" => DATA <= x"4C";
      when x"997" => DATA <= x"A4";
      when x"998" => DATA <= x"DA";
      when x"999" => DATA <= x"B0";
      when x"99A" => DATA <= x"2D";
      when x"99B" => DATA <= x"38";
      when x"99C" => DATA <= x"A5";
      when x"99D" => DATA <= x"66";
      when x"99E" => DATA <= x"E5";
      when x"99F" => DATA <= x"5E";
      when x"9A0" => DATA <= x"85";
      when x"9A1" => DATA <= x"5E";
      when x"9A2" => DATA <= x"A5";
      when x"9A3" => DATA <= x"65";
      when x"9A4" => DATA <= x"E5";
      when x"9A5" => DATA <= x"5D";
      when x"9A6" => DATA <= x"85";
      when x"9A7" => DATA <= x"5D";
      when x"9A8" => DATA <= x"A5";
      when x"9A9" => DATA <= x"64";
      when x"9AA" => DATA <= x"E5";
      when x"9AB" => DATA <= x"5C";
      when x"9AC" => DATA <= x"85";
      when x"9AD" => DATA <= x"5C";
      when x"9AE" => DATA <= x"A5";
      when x"9AF" => DATA <= x"63";
      when x"9B0" => DATA <= x"E5";
      when x"9B1" => DATA <= x"5B";
      when x"9B2" => DATA <= x"85";
      when x"9B3" => DATA <= x"5B";
      when x"9B4" => DATA <= x"A5";
      when x"9B5" => DATA <= x"62";
      when x"9B6" => DATA <= x"E5";
      when x"9B7" => DATA <= x"5A";
      when x"9B8" => DATA <= x"85";
      when x"9B9" => DATA <= x"5A";
      when x"9BA" => DATA <= x"A5";
      when x"9BB" => DATA <= x"5F";
      when x"9BC" => DATA <= x"85";
      when x"9BD" => DATA <= x"57";
      when x"9BE" => DATA <= x"4C";
      when x"9BF" => DATA <= x"98";
      when x"9C0" => DATA <= x"DA";
      when x"9C1" => DATA <= x"18";
      when x"9C2" => DATA <= x"20";
      when x"9C3" => DATA <= x"B4";
      when x"9C4" => DATA <= x"D6";
      when x"9C5" => DATA <= x"4C";
      when x"9C6" => DATA <= x"9B";
      when x"9C7" => DATA <= x"DA";
      when x"9C8" => DATA <= x"38";
      when x"9C9" => DATA <= x"A5";
      when x"9CA" => DATA <= x"5E";
      when x"9CB" => DATA <= x"E5";
      when x"9CC" => DATA <= x"66";
      when x"9CD" => DATA <= x"85";
      when x"9CE" => DATA <= x"5E";
      when x"9CF" => DATA <= x"A5";
      when x"9D0" => DATA <= x"5D";
      when x"9D1" => DATA <= x"E5";
      when x"9D2" => DATA <= x"65";
      when x"9D3" => DATA <= x"85";
      when x"9D4" => DATA <= x"5D";
      when x"9D5" => DATA <= x"A5";
      when x"9D6" => DATA <= x"5C";
      when x"9D7" => DATA <= x"E5";
      when x"9D8" => DATA <= x"64";
      when x"9D9" => DATA <= x"85";
      when x"9DA" => DATA <= x"5C";
      when x"9DB" => DATA <= x"A5";
      when x"9DC" => DATA <= x"5B";
      when x"9DD" => DATA <= x"E5";
      when x"9DE" => DATA <= x"63";
      when x"9DF" => DATA <= x"85";
      when x"9E0" => DATA <= x"5B";
      when x"9E1" => DATA <= x"A5";
      when x"9E2" => DATA <= x"5A";
      when x"9E3" => DATA <= x"E5";
      when x"9E4" => DATA <= x"62";
      when x"9E5" => DATA <= x"85";
      when x"9E6" => DATA <= x"5A";
      when x"9E7" => DATA <= x"4C";
      when x"9E8" => DATA <= x"98";
      when x"9E9" => DATA <= x"DA";
      when x"9EA" => DATA <= x"00";
      when x"9EB" => DATA <= x"20";
      when x"9EC" => DATA <= x"FC";
      when x"9ED" => DATA <= x"D0";
      when x"9EE" => DATA <= x"A9";
      when x"9EF" => DATA <= x"C7";
      when x"9F0" => DATA <= x"48";
      when x"9F1" => DATA <= x"A2";
      when x"9F2" => DATA <= x"C8";
      when x"9F3" => DATA <= x"4C";
      when x"9F4" => DATA <= x"0B";
      when x"9F5" => DATA <= x"D1";
      when x"9F6" => DATA <= x"A9";
      when x"9F7" => DATA <= x"5D";
      when x"9F8" => DATA <= x"D0";
      when x"9F9" => DATA <= x"12";
      when x"9FA" => DATA <= x"A9";
      when x"9FB" => DATA <= x"66";
      when x"9FC" => DATA <= x"D0";
      when x"9FD" => DATA <= x"0E";
      when x"9FE" => DATA <= x"A9";
      when x"9FF" => DATA <= x"6F";
      when x"A00" => DATA <= x"D0";
      when x"A01" => DATA <= x"0A";
      when x"A02" => DATA <= x"A9";
      when x"A03" => DATA <= x"76";
      when x"A04" => DATA <= x"D0";
      when x"A05" => DATA <= x"06";
      when x"A06" => DATA <= x"A9";
      when x"A07" => DATA <= x"7D";
      when x"A08" => DATA <= x"D0";
      when x"A09" => DATA <= x"02";
      when x"A0A" => DATA <= x"A9";
      when x"A0B" => DATA <= x"84";
      when x"A0C" => DATA <= x"48";
      when x"A0D" => DATA <= x"20";
      when x"A0E" => DATA <= x"5D";
      when x"A0F" => DATA <= x"D8";
      when x"A10" => DATA <= x"20";
      when x"A11" => DATA <= x"FC";
      when x"A12" => DATA <= x"D0";
      when x"A13" => DATA <= x"20";
      when x"A14" => DATA <= x"70";
      when x"A15" => DATA <= x"D8";
      when x"A16" => DATA <= x"E6";
      when x"A17" => DATA <= x"04";
      when x"A18" => DATA <= x"20";
      when x"A19" => DATA <= x"04";
      when x"A1A" => DATA <= x"D8";
      when x"A1B" => DATA <= x"A5";
      when x"A1C" => DATA <= x"5F";
      when x"A1D" => DATA <= x"29";
      when x"A1E" => DATA <= x"80";
      when x"A1F" => DATA <= x"85";
      when x"A20" => DATA <= x"5F";
      when x"A21" => DATA <= x"A0";
      when x"A22" => DATA <= x"00";
      when x"A23" => DATA <= x"A5";
      when x"A24" => DATA <= x"57";
      when x"A25" => DATA <= x"29";
      when x"A26" => DATA <= x"80";
      when x"A27" => DATA <= x"C5";
      when x"A28" => DATA <= x"5F";
      when x"A29" => DATA <= x"D0";
      when x"A2A" => DATA <= x"0D";
      when x"A2B" => DATA <= x"A2";
      when x"A2C" => DATA <= x"00";
      when x"A2D" => DATA <= x"B5";
      when x"A2E" => DATA <= x"61";
      when x"A2F" => DATA <= x"D5";
      when x"A30" => DATA <= x"59";
      when x"A31" => DATA <= x"D0";
      when x"A32" => DATA <= x"0A";
      when x"A33" => DATA <= x"E8";
      when x"A34" => DATA <= x"E0";
      when x"A35" => DATA <= x"05";
      when x"A36" => DATA <= x"D0";
      when x"A37" => DATA <= x"F5";
      when x"A38" => DATA <= x"08";
      when x"A39" => DATA <= x"A6";
      when x"A3A" => DATA <= x"04";
      when x"A3B" => DATA <= x"28";
      when x"A3C" => DATA <= x"60";
      when x"A3D" => DATA <= x"6A";
      when x"A3E" => DATA <= x"45";
      when x"A3F" => DATA <= x"5F";
      when x"A40" => DATA <= x"2A";
      when x"A41" => DATA <= x"A9";
      when x"A42" => DATA <= x"01";
      when x"A43" => DATA <= x"D0";
      when x"A44" => DATA <= x"F3";
      when x"A45" => DATA <= x"20";
      when x"A46" => DATA <= x"86";
      when x"A47" => DATA <= x"D6";
      when x"A48" => DATA <= x"F0";
      when x"A49" => DATA <= x"F2";
      when x"A4A" => DATA <= x"20";
      when x"A4B" => DATA <= x"04";
      when x"A4C" => DATA <= x"D8";
      when x"A4D" => DATA <= x"D0";
      when x"A4E" => DATA <= x"03";
      when x"A4F" => DATA <= x"4C";
      when x"A50" => DATA <= x"A4";
      when x"A51" => DATA <= x"DA";
      when x"A52" => DATA <= x"18";
      when x"A53" => DATA <= x"A5";
      when x"A54" => DATA <= x"59";
      when x"A55" => DATA <= x"65";
      when x"A56" => DATA <= x"61";
      when x"A57" => DATA <= x"85";
      when x"A58" => DATA <= x"59";
      when x"A59" => DATA <= x"90";
      when x"A5A" => DATA <= x"02";
      when x"A5B" => DATA <= x"E6";
      when x"A5C" => DATA <= x"58";
      when x"A5D" => DATA <= x"38";
      when x"A5E" => DATA <= x"A5";
      when x"A5F" => DATA <= x"59";
      when x"A60" => DATA <= x"E9";
      when x"A61" => DATA <= x"80";
      when x"A62" => DATA <= x"85";
      when x"A63" => DATA <= x"59";
      when x"A64" => DATA <= x"B0";
      when x"A65" => DATA <= x"02";
      when x"A66" => DATA <= x"C6";
      when x"A67" => DATA <= x"58";
      when x"A68" => DATA <= x"A2";
      when x"A69" => DATA <= x"05";
      when x"A6A" => DATA <= x"A0";
      when x"A6B" => DATA <= x"00";
      when x"A6C" => DATA <= x"B5";
      when x"A6D" => DATA <= x"59";
      when x"A6E" => DATA <= x"95";
      when x"A6F" => DATA <= x"66";
      when x"A70" => DATA <= x"94";
      when x"A71" => DATA <= x"59";
      when x"A72" => DATA <= x"CA";
      when x"A73" => DATA <= x"D0";
      when x"A74" => DATA <= x"F7";
      when x"A75" => DATA <= x"A5";
      when x"A76" => DATA <= x"57";
      when x"A77" => DATA <= x"45";
      when x"A78" => DATA <= x"5F";
      when x"A79" => DATA <= x"85";
      when x"A7A" => DATA <= x"57";
      when x"A7B" => DATA <= x"A0";
      when x"A7C" => DATA <= x"20";
      when x"A7D" => DATA <= x"20";
      when x"A7E" => DATA <= x"FB";
      when x"A7F" => DATA <= x"D6";
      when x"A80" => DATA <= x"A5";
      when x"A81" => DATA <= x"67";
      when x"A82" => DATA <= x"10";
      when x"A83" => DATA <= x"04";
      when x"A84" => DATA <= x"18";
      when x"A85" => DATA <= x"20";
      when x"A86" => DATA <= x"42";
      when x"A87" => DATA <= x"D6";
      when x"A88" => DATA <= x"20";
      when x"A89" => DATA <= x"FB";
      when x"A8A" => DATA <= x"D6";
      when x"A8B" => DATA <= x"06";
      when x"A8C" => DATA <= x"6B";
      when x"A8D" => DATA <= x"26";
      when x"A8E" => DATA <= x"6A";
      when x"A8F" => DATA <= x"26";
      when x"A90" => DATA <= x"69";
      when x"A91" => DATA <= x"26";
      when x"A92" => DATA <= x"68";
      when x"A93" => DATA <= x"26";
      when x"A94" => DATA <= x"67";
      when x"A95" => DATA <= x"88";
      when x"A96" => DATA <= x"D0";
      when x"A97" => DATA <= x"E8";
      when x"A98" => DATA <= x"20";
      when x"A99" => DATA <= x"C8";
      when x"A9A" => DATA <= x"D7";
      when x"A9B" => DATA <= x"20";
      when x"A9C" => DATA <= x"80";
      when x"A9D" => DATA <= x"D8";
      when x"A9E" => DATA <= x"A5";
      when x"A9F" => DATA <= x"58";
      when x"AA0" => DATA <= x"F0";
      when x"AA1" => DATA <= x"0B";
      when x"AA2" => DATA <= x"10";
      when x"AA3" => DATA <= x"03";
      when x"AA4" => DATA <= x"A2";
      when x"AA5" => DATA <= x"08";
      when x"AA6" => DATA <= x"A9";
      when x"AA7" => DATA <= x"00";
      when x"AA8" => DATA <= x"95";
      when x"AA9" => DATA <= x"56";
      when x"AAA" => DATA <= x"CA";
      when x"AAB" => DATA <= x"D0";
      when x"AAC" => DATA <= x"FB";
      when x"AAD" => DATA <= x"60";
      when x"AAE" => DATA <= x"20";
      when x"AAF" => DATA <= x"31";
      when x"AB0" => DATA <= x"D8";
      when x"AB1" => DATA <= x"20";
      when x"AB2" => DATA <= x"8D";
      when x"AB3" => DATA <= x"DE";
      when x"AB4" => DATA <= x"D0";
      when x"AB5" => DATA <= x"26";
      when x"AB6" => DATA <= x"20";
      when x"AB7" => DATA <= x"86";
      when x"AB8" => DATA <= x"D6";
      when x"AB9" => DATA <= x"F0";
      when x"ABA" => DATA <= x"EC";
      when x"ABB" => DATA <= x"20";
      when x"ABC" => DATA <= x"C3";
      when x"ABD" => DATA <= x"D6";
      when x"ABE" => DATA <= x"20";
      when x"ABF" => DATA <= x"E5";
      when x"AC0" => DATA <= x"D1";
      when x"AC1" => DATA <= x"D0";
      when x"AC2" => DATA <= x"23";
      when x"AC3" => DATA <= x"60";
      when x"AC4" => DATA <= x"20";
      when x"AC5" => DATA <= x"EB";
      when x"AC6" => DATA <= x"D0";
      when x"AC7" => DATA <= x"20";
      when x"AC8" => DATA <= x"9E";
      when x"AC9" => DATA <= x"DB";
      when x"ACA" => DATA <= x"20";
      when x"ACB" => DATA <= x"3D";
      when x"ACC" => DATA <= x"D8";
      when x"ACD" => DATA <= x"20";
      when x"ACE" => DATA <= x"E6";
      when x"ACF" => DATA <= x"DC";
      when x"AD0" => DATA <= x"20";
      when x"AD1" => DATA <= x"9E";
      when x"AD2" => DATA <= x"DB";
      when x"AD3" => DATA <= x"20";
      when x"AD4" => DATA <= x"23";
      when x"AD5" => DATA <= x"D9";
      when x"AD6" => DATA <= x"20";
      when x"AD7" => DATA <= x"F1";
      when x"AD8" => DATA <= x"DC";
      when x"AD9" => DATA <= x"20";
      when x"ADA" => DATA <= x"9E";
      when x"ADB" => DATA <= x"DB";
      when x"ADC" => DATA <= x"20";
      when x"ADD" => DATA <= x"86";
      when x"ADE" => DATA <= x"D6";
      when x"ADF" => DATA <= x"F0";
      when x"AE0" => DATA <= x"CC";
      when x"AE1" => DATA <= x"20";
      when x"AE2" => DATA <= x"04";
      when x"AE3" => DATA <= x"D8";
      when x"AE4" => DATA <= x"F0";
      when x"AE5" => DATA <= x"C1";
      when x"AE6" => DATA <= x"A5";
      when x"AE7" => DATA <= x"57";
      when x"AE8" => DATA <= x"45";
      when x"AE9" => DATA <= x"5F";
      when x"AEA" => DATA <= x"85";
      when x"AEB" => DATA <= x"57";
      when x"AEC" => DATA <= x"38";
      when x"AED" => DATA <= x"A5";
      when x"AEE" => DATA <= x"59";
      when x"AEF" => DATA <= x"E5";
      when x"AF0" => DATA <= x"61";
      when x"AF1" => DATA <= x"85";
      when x"AF2" => DATA <= x"59";
      when x"AF3" => DATA <= x"B0";
      when x"AF4" => DATA <= x"02";
      when x"AF5" => DATA <= x"C6";
      when x"AF6" => DATA <= x"58";
      when x"AF7" => DATA <= x"18";
      when x"AF8" => DATA <= x"A5";
      when x"AF9" => DATA <= x"59";
      when x"AFA" => DATA <= x"69";
      when x"AFB" => DATA <= x"81";
      when x"AFC" => DATA <= x"85";
      when x"AFD" => DATA <= x"59";
      when x"AFE" => DATA <= x"90";
      when x"AFF" => DATA <= x"02";
      when x"B00" => DATA <= x"E6";
      when x"B01" => DATA <= x"58";
      when x"B02" => DATA <= x"A2";
      when x"B03" => DATA <= x"05";
      when x"B04" => DATA <= x"B5";
      when x"B05" => DATA <= x"59";
      when x"B06" => DATA <= x"95";
      when x"B07" => DATA <= x"66";
      when x"B08" => DATA <= x"CA";
      when x"B09" => DATA <= x"D0";
      when x"B0A" => DATA <= x"F9";
      when x"B0B" => DATA <= x"46";
      when x"B0C" => DATA <= x"67";
      when x"B0D" => DATA <= x"66";
      when x"B0E" => DATA <= x"68";
      when x"B0F" => DATA <= x"66";
      when x"B10" => DATA <= x"69";
      when x"B11" => DATA <= x"66";
      when x"B12" => DATA <= x"6A";
      when x"B13" => DATA <= x"66";
      when x"B14" => DATA <= x"6B";
      when x"B15" => DATA <= x"20";
      when x"B16" => DATA <= x"FB";
      when x"B17" => DATA <= x"D6";
      when x"B18" => DATA <= x"A2";
      when x"B19" => DATA <= x"27";
      when x"B1A" => DATA <= x"A5";
      when x"B1B" => DATA <= x"67";
      when x"B1C" => DATA <= x"C5";
      when x"B1D" => DATA <= x"62";
      when x"B1E" => DATA <= x"D0";
      when x"B1F" => DATA <= x"16";
      when x"B20" => DATA <= x"A5";
      when x"B21" => DATA <= x"68";
      when x"B22" => DATA <= x"C5";
      when x"B23" => DATA <= x"63";
      when x"B24" => DATA <= x"D0";
      when x"B25" => DATA <= x"10";
      when x"B26" => DATA <= x"A5";
      when x"B27" => DATA <= x"69";
      when x"B28" => DATA <= x"C5";
      when x"B29" => DATA <= x"64";
      when x"B2A" => DATA <= x"D0";
      when x"B2B" => DATA <= x"0A";
      when x"B2C" => DATA <= x"A5";
      when x"B2D" => DATA <= x"6A";
      when x"B2E" => DATA <= x"C5";
      when x"B2F" => DATA <= x"65";
      when x"B30" => DATA <= x"D0";
      when x"B31" => DATA <= x"04";
      when x"B32" => DATA <= x"A5";
      when x"B33" => DATA <= x"6B";
      when x"B34" => DATA <= x"C5";
      when x"B35" => DATA <= x"66";
      when x"B36" => DATA <= x"90";
      when x"B37" => DATA <= x"24";
      when x"B38" => DATA <= x"A5";
      when x"B39" => DATA <= x"6B";
      when x"B3A" => DATA <= x"E5";
      when x"B3B" => DATA <= x"66";
      when x"B3C" => DATA <= x"85";
      when x"B3D" => DATA <= x"6B";
      when x"B3E" => DATA <= x"A5";
      when x"B3F" => DATA <= x"6A";
      when x"B40" => DATA <= x"E5";
      when x"B41" => DATA <= x"65";
      when x"B42" => DATA <= x"85";
      when x"B43" => DATA <= x"6A";
      when x"B44" => DATA <= x"A5";
      when x"B45" => DATA <= x"69";
      when x"B46" => DATA <= x"E5";
      when x"B47" => DATA <= x"64";
      when x"B48" => DATA <= x"85";
      when x"B49" => DATA <= x"69";
      when x"B4A" => DATA <= x"A5";
      when x"B4B" => DATA <= x"68";
      when x"B4C" => DATA <= x"E5";
      when x"B4D" => DATA <= x"63";
      when x"B4E" => DATA <= x"85";
      when x"B4F" => DATA <= x"68";
      when x"B50" => DATA <= x"A5";
      when x"B51" => DATA <= x"67";
      when x"B52" => DATA <= x"E5";
      when x"B53" => DATA <= x"62";
      when x"B54" => DATA <= x"85";
      when x"B55" => DATA <= x"67";
      when x"B56" => DATA <= x"A5";
      when x"B57" => DATA <= x"5E";
      when x"B58" => DATA <= x"09";
      when x"B59" => DATA <= x"01";
      when x"B5A" => DATA <= x"85";
      when x"B5B" => DATA <= x"5E";
      when x"B5C" => DATA <= x"20";
      when x"B5D" => DATA <= x"CD";
      when x"B5E" => DATA <= x"D6";
      when x"B5F" => DATA <= x"06";
      when x"B60" => DATA <= x"6B";
      when x"B61" => DATA <= x"26";
      when x"B62" => DATA <= x"6A";
      when x"B63" => DATA <= x"26";
      when x"B64" => DATA <= x"69";
      when x"B65" => DATA <= x"26";
      when x"B66" => DATA <= x"68";
      when x"B67" => DATA <= x"26";
      when x"B68" => DATA <= x"67";
      when x"B69" => DATA <= x"CA";
      when x"B6A" => DATA <= x"D0";
      when x"B6B" => DATA <= x"AE";
      when x"B6C" => DATA <= x"4C";
      when x"B6D" => DATA <= x"98";
      when x"B6E" => DATA <= x"DA";
      when x"B6F" => DATA <= x"20";
      when x"B70" => DATA <= x"EB";
      when x"B71" => DATA <= x"D0";
      when x"B72" => DATA <= x"20";
      when x"B73" => DATA <= x"86";
      when x"B74" => DATA <= x"D6";
      when x"B75" => DATA <= x"F0";
      when x"B76" => DATA <= x"26";
      when x"B77" => DATA <= x"10";
      when x"B78" => DATA <= x"01";
      when x"B79" => DATA <= x"00";
      when x"B7A" => DATA <= x"20";
      when x"B7B" => DATA <= x"31";
      when x"B7C" => DATA <= x"D8";
      when x"B7D" => DATA <= x"A5";
      when x"B7E" => DATA <= x"59";
      when x"B7F" => DATA <= x"4A";
      when x"B80" => DATA <= x"69";
      when x"B81" => DATA <= x"40";
      when x"B82" => DATA <= x"85";
      when x"B83" => DATA <= x"59";
      when x"B84" => DATA <= x"A9";
      when x"B85" => DATA <= x"05";
      when x"B86" => DATA <= x"85";
      when x"B87" => DATA <= x"6E";
      when x"B88" => DATA <= x"20";
      when x"B89" => DATA <= x"27";
      when x"B8A" => DATA <= x"D8";
      when x"B8B" => DATA <= x"20";
      when x"B8C" => DATA <= x"AA";
      when x"B8D" => DATA <= x"DB";
      when x"B8E" => DATA <= x"20";
      when x"B8F" => DATA <= x"B6";
      when x"B90" => DATA <= x"DA";
      when x"B91" => DATA <= x"20";
      when x"B92" => DATA <= x"A2";
      when x"B93" => DATA <= x"DB";
      when x"B94" => DATA <= x"20";
      when x"B95" => DATA <= x"3C";
      when x"B96" => DATA <= x"D9";
      when x"B97" => DATA <= x"C6";
      when x"B98" => DATA <= x"59";
      when x"B99" => DATA <= x"C6";
      when x"B9A" => DATA <= x"6E";
      when x"B9B" => DATA <= x"D0";
      when x"B9C" => DATA <= x"EB";
      when x"B9D" => DATA <= x"60";
      when x"B9E" => DATA <= x"A9";
      when x"B9F" => DATA <= x"D4";
      when x"BA0" => DATA <= x"D0";
      when x"BA1" => DATA <= x"0A";
      when x"BA2" => DATA <= x"A9";
      when x"BA3" => DATA <= x"CA";
      when x"BA4" => DATA <= x"D0";
      when x"BA5" => DATA <= x"06";
      when x"BA6" => DATA <= x"A9";
      when x"BA7" => DATA <= x"CF";
      when x"BA8" => DATA <= x"D0";
      when x"BA9" => DATA <= x"02";
      when x"BAA" => DATA <= x"A9";
      when x"BAB" => DATA <= x"C5";
      when x"BAC" => DATA <= x"85";
      when x"BAD" => DATA <= x"6F";
      when x"BAE" => DATA <= x"A9";
      when x"BAF" => DATA <= x"03";
      when x"BB0" => DATA <= x"85";
      when x"BB1" => DATA <= x"70";
      when x"BB2" => DATA <= x"60";
      when x"BB3" => DATA <= x"20";
      when x"BB4" => DATA <= x"EB";
      when x"BB5" => DATA <= x"D0";
      when x"BB6" => DATA <= x"20";
      when x"BB7" => DATA <= x"86";
      when x"BB8" => DATA <= x"D6";
      when x"BB9" => DATA <= x"F0";
      when x"BBA" => DATA <= x"02";
      when x"BBB" => DATA <= x"10";
      when x"BBC" => DATA <= x"01";
      when x"BBD" => DATA <= x"00";
      when x"BBE" => DATA <= x"A5";
      when x"BBF" => DATA <= x"59";
      when x"BC0" => DATA <= x"48";
      when x"BC1" => DATA <= x"A9";
      when x"BC2" => DATA <= x"81";
      when x"BC3" => DATA <= x"85";
      when x"BC4" => DATA <= x"59";
      when x"BC5" => DATA <= x"20";
      when x"BC6" => DATA <= x"C7";
      when x"BC7" => DATA <= x"D8";
      when x"BC8" => DATA <= x"A9";
      when x"BC9" => DATA <= x"C0";
      when x"BCA" => DATA <= x"85";
      when x"BCB" => DATA <= x"62";
      when x"BCC" => DATA <= x"A9";
      when x"BCD" => DATA <= x"81";
      when x"BCE" => DATA <= x"85";
      when x"BCF" => DATA <= x"61";
      when x"BD0" => DATA <= x"85";
      when x"BD1" => DATA <= x"5F";
      when x"BD2" => DATA <= x"20";
      when x"BD3" => DATA <= x"41";
      when x"BD4" => DATA <= x"D9";
      when x"BD5" => DATA <= x"E6";
      when x"BD6" => DATA <= x"59";
      when x"BD7" => DATA <= x"A9";
      when x"BD8" => DATA <= x"FE";
      when x"BD9" => DATA <= x"A0";
      when x"BDA" => DATA <= x"DB";
      when x"BDB" => DATA <= x"20";
      when x"BDC" => DATA <= x"27";
      when x"BDD" => DATA <= x"DC";
      when x"BDE" => DATA <= x"20";
      when x"BDF" => DATA <= x"31";
      when x"BE0" => DATA <= x"D8";
      when x"BE1" => DATA <= x"68";
      when x"BE2" => DATA <= x"38";
      when x"BE3" => DATA <= x"E9";
      when x"BE4" => DATA <= x"81";
      when x"BE5" => DATA <= x"20";
      when x"BE6" => DATA <= x"B2";
      when x"BE7" => DATA <= x"D7";
      when x"BE8" => DATA <= x"A9";
      when x"BE9" => DATA <= x"F9";
      when x"BEA" => DATA <= x"85";
      when x"BEB" => DATA <= x"6F";
      when x"BEC" => DATA <= x"A9";
      when x"BED" => DATA <= x"DB";
      when x"BEE" => DATA <= x"85";
      when x"BEF" => DATA <= x"70";
      when x"BF0" => DATA <= x"20";
      when x"BF1" => DATA <= x"45";
      when x"BF2" => DATA <= x"DA";
      when x"BF3" => DATA <= x"20";
      when x"BF4" => DATA <= x"AA";
      when x"BF5" => DATA <= x"DB";
      when x"BF6" => DATA <= x"4C";
      when x"BF7" => DATA <= x"3C";
      when x"BF8" => DATA <= x"D9";
      when x"BF9" => DATA <= x"80";
      when x"BFA" => DATA <= x"31";
      when x"BFB" => DATA <= x"72";
      when x"BFC" => DATA <= x"17";
      when x"BFD" => DATA <= x"F8";
      when x"BFE" => DATA <= x"07";
      when x"BFF" => DATA <= x"85";
      when x"C00" => DATA <= x"17";
      when x"C01" => DATA <= x"6E";
      when x"C02" => DATA <= x"D4";
      when x"C03" => DATA <= x"85";
      when x"C04" => DATA <= x"80";
      when x"C05" => DATA <= x"28";
      when x"C06" => DATA <= x"C7";
      when x"C07" => DATA <= x"12";
      when x"C08" => DATA <= x"A0";
      when x"C09" => DATA <= x"84";
      when x"C0A" => DATA <= x"70";
      when x"C0B" => DATA <= x"4E";
      when x"C0C" => DATA <= x"5F";
      when x"C0D" => DATA <= x"F2";
      when x"C0E" => DATA <= x"81";
      when x"C0F" => DATA <= x"00";
      when x"C10" => DATA <= x"00";
      when x"C11" => DATA <= x"FE";
      when x"C12" => DATA <= x"EF";
      when x"C13" => DATA <= x"84";
      when x"C14" => DATA <= x"0F";
      when x"C15" => DATA <= x"FF";
      when x"C16" => DATA <= x"DA";
      when x"C17" => DATA <= x"E1";
      when x"C18" => DATA <= x"81";
      when x"C19" => DATA <= x"7F";
      when x"C1A" => DATA <= x"FF";
      when x"C1B" => DATA <= x"FF";
      when x"C1C" => DATA <= x"93";
      when x"C1D" => DATA <= x"82";
      when x"C1E" => DATA <= x"40";
      when x"C1F" => DATA <= x"00";
      when x"C20" => DATA <= x"00";
      when x"C21" => DATA <= x"0C";
      when x"C22" => DATA <= x"7F";
      when x"C23" => DATA <= x"4F";
      when x"C24" => DATA <= x"99";
      when x"C25" => DATA <= x"1F";
      when x"C26" => DATA <= x"65";
      when x"C27" => DATA <= x"85";
      when x"C28" => DATA <= x"71";
      when x"C29" => DATA <= x"84";
      when x"C2A" => DATA <= x"72";
      when x"C2B" => DATA <= x"20";
      when x"C2C" => DATA <= x"31";
      when x"C2D" => DATA <= x"D8";
      when x"C2E" => DATA <= x"A0";
      when x"C2F" => DATA <= x"00";
      when x"C30" => DATA <= x"B1";
      when x"C31" => DATA <= x"71";
      when x"C32" => DATA <= x"85";
      when x"C33" => DATA <= x"6C";
      when x"C34" => DATA <= x"E6";
      when x"C35" => DATA <= x"71";
      when x"C36" => DATA <= x"D0";
      when x"C37" => DATA <= x"02";
      when x"C38" => DATA <= x"E6";
      when x"C39" => DATA <= x"72";
      when x"C3A" => DATA <= x"A5";
      when x"C3B" => DATA <= x"71";
      when x"C3C" => DATA <= x"85";
      when x"C3D" => DATA <= x"6F";
      when x"C3E" => DATA <= x"A5";
      when x"C3F" => DATA <= x"72";
      when x"C40" => DATA <= x"85";
      when x"C41" => DATA <= x"70";
      when x"C42" => DATA <= x"20";
      when x"C43" => DATA <= x"E5";
      when x"C44" => DATA <= x"D1";
      when x"C45" => DATA <= x"20";
      when x"C46" => DATA <= x"AA";
      when x"C47" => DATA <= x"DB";
      when x"C48" => DATA <= x"20";
      when x"C49" => DATA <= x"B6";
      when x"C4A" => DATA <= x"DA";
      when x"C4B" => DATA <= x"18";
      when x"C4C" => DATA <= x"A5";
      when x"C4D" => DATA <= x"71";
      when x"C4E" => DATA <= x"69";
      when x"C4F" => DATA <= x"05";
      when x"C50" => DATA <= x"85";
      when x"C51" => DATA <= x"71";
      when x"C52" => DATA <= x"85";
      when x"C53" => DATA <= x"6F";
      when x"C54" => DATA <= x"A5";
      when x"C55" => DATA <= x"72";
      when x"C56" => DATA <= x"69";
      when x"C57" => DATA <= x"00";
      when x"C58" => DATA <= x"85";
      when x"C59" => DATA <= x"72";
      when x"C5A" => DATA <= x"85";
      when x"C5B" => DATA <= x"70";
      when x"C5C" => DATA <= x"20";
      when x"C5D" => DATA <= x"3C";
      when x"C5E" => DATA <= x"D9";
      when x"C5F" => DATA <= x"C6";
      when x"C60" => DATA <= x"6C";
      when x"C61" => DATA <= x"D0";
      when x"C62" => DATA <= x"E2";
      when x"C63" => DATA <= x"60";
      when x"C64" => DATA <= x"20";
      when x"C65" => DATA <= x"EB";
      when x"C66" => DATA <= x"D0";
      when x"C67" => DATA <= x"20";
      when x"C68" => DATA <= x"86";
      when x"C69" => DATA <= x"D6";
      when x"C6A" => DATA <= x"F0";
      when x"C6B" => DATA <= x"0D";
      when x"C6C" => DATA <= x"10";
      when x"C6D" => DATA <= x"0C";
      when x"C6E" => DATA <= x"A9";
      when x"C6F" => DATA <= x"00";
      when x"C70" => DATA <= x"85";
      when x"C71" => DATA <= x"57";
      when x"C72" => DATA <= x"20";
      when x"C73" => DATA <= x"7A";
      when x"C74" => DATA <= x"DC";
      when x"C75" => DATA <= x"A9";
      when x"C76" => DATA <= x"80";
      when x"C77" => DATA <= x"85";
      when x"C78" => DATA <= x"57";
      when x"C79" => DATA <= x"60";
      when x"C7A" => DATA <= x"A5";
      when x"C7B" => DATA <= x"59";
      when x"C7C" => DATA <= x"C9";
      when x"C7D" => DATA <= x"81";
      when x"C7E" => DATA <= x"90";
      when x"C7F" => DATA <= x"0C";
      when x"C80" => DATA <= x"20";
      when x"C81" => DATA <= x"AE";
      when x"C82" => DATA <= x"DA";
      when x"C83" => DATA <= x"20";
      when x"C84" => DATA <= x"8C";
      when x"C85" => DATA <= x"DC";
      when x"C86" => DATA <= x"20";
      when x"C87" => DATA <= x"93";
      when x"C88" => DATA <= x"DD";
      when x"C89" => DATA <= x"4C";
      when x"C8A" => DATA <= x"39";
      when x"C8B" => DATA <= x"D9";
      when x"C8C" => DATA <= x"A5";
      when x"C8D" => DATA <= x"59";
      when x"C8E" => DATA <= x"C9";
      when x"C8F" => DATA <= x"73";
      when x"C90" => DATA <= x"90";
      when x"C91" => DATA <= x"E7";
      when x"C92" => DATA <= x"20";
      when x"C93" => DATA <= x"2C";
      when x"C94" => DATA <= x"D8";
      when x"C95" => DATA <= x"20";
      when x"C96" => DATA <= x"C7";
      when x"C97" => DATA <= x"D8";
      when x"C98" => DATA <= x"A9";
      when x"C99" => DATA <= x"80";
      when x"C9A" => DATA <= x"85";
      when x"C9B" => DATA <= x"61";
      when x"C9C" => DATA <= x"85";
      when x"C9D" => DATA <= x"62";
      when x"C9E" => DATA <= x"85";
      when x"C9F" => DATA <= x"5F";
      when x"CA0" => DATA <= x"20";
      when x"CA1" => DATA <= x"41";
      when x"CA2" => DATA <= x"D9";
      when x"CA3" => DATA <= x"A9";
      when x"CA4" => DATA <= x"B0";
      when x"CA5" => DATA <= x"A0";
      when x"CA6" => DATA <= x"DC";
      when x"CA7" => DATA <= x"20";
      when x"CA8" => DATA <= x"27";
      when x"CA9" => DATA <= x"DC";
      when x"CAA" => DATA <= x"20";
      when x"CAB" => DATA <= x"A6";
      when x"CAC" => DATA <= x"DB";
      when x"CAD" => DATA <= x"4C";
      when x"CAE" => DATA <= x"45";
      when x"CAF" => DATA <= x"DA";
      when x"CB0" => DATA <= x"09";
      when x"CB1" => DATA <= x"85";
      when x"CB2" => DATA <= x"A3";
      when x"CB3" => DATA <= x"59";
      when x"CB4" => DATA <= x"E8";
      when x"CB5" => DATA <= x"67";
      when x"CB6" => DATA <= x"80";
      when x"CB7" => DATA <= x"1C";
      when x"CB8" => DATA <= x"9D";
      when x"CB9" => DATA <= x"07";
      when x"CBA" => DATA <= x"36";
      when x"CBB" => DATA <= x"80";
      when x"CBC" => DATA <= x"57";
      when x"CBD" => DATA <= x"BB";
      when x"CBE" => DATA <= x"78";
      when x"CBF" => DATA <= x"DF";
      when x"CC0" => DATA <= x"80";
      when x"CC1" => DATA <= x"CA";
      when x"CC2" => DATA <= x"9A";
      when x"CC3" => DATA <= x"0E";
      when x"CC4" => DATA <= x"83";
      when x"CC5" => DATA <= x"84";
      when x"CC6" => DATA <= x"8C";
      when x"CC7" => DATA <= x"BB";
      when x"CC8" => DATA <= x"CA";
      when x"CC9" => DATA <= x"6E";
      when x"CCA" => DATA <= x"81";
      when x"CCB" => DATA <= x"95";
      when x"CCC" => DATA <= x"96";
      when x"CCD" => DATA <= x"06";
      when x"CCE" => DATA <= x"DE";
      when x"CCF" => DATA <= x"81";
      when x"CD0" => DATA <= x"0A";
      when x"CD1" => DATA <= x"C7";
      when x"CD2" => DATA <= x"6C";
      when x"CD3" => DATA <= x"52";
      when x"CD4" => DATA <= x"7F";
      when x"CD5" => DATA <= x"7D";
      when x"CD6" => DATA <= x"AD";
      when x"CD7" => DATA <= x"90";
      when x"CD8" => DATA <= x"A1";
      when x"CD9" => DATA <= x"82";
      when x"CDA" => DATA <= x"FB";
      when x"CDB" => DATA <= x"62";
      when x"CDC" => DATA <= x"57";
      when x"CDD" => DATA <= x"2F";
      when x"CDE" => DATA <= x"80";
      when x"CDF" => DATA <= x"6D";
      when x"CE0" => DATA <= x"63";
      when x"CE1" => DATA <= x"38";
      when x"CE2" => DATA <= x"2C";
      when x"CE3" => DATA <= x"20";
      when x"CE4" => DATA <= x"EB";
      when x"CE5" => DATA <= x"D0";
      when x"CE6" => DATA <= x"20";
      when x"CE7" => DATA <= x"24";
      when x"CE8" => DATA <= x"DD";
      when x"CE9" => DATA <= x"E6";
      when x"CEA" => DATA <= x"6E";
      when x"CEB" => DATA <= x"4C";
      when x"CEC" => DATA <= x"F4";
      when x"CED" => DATA <= x"DC";
      when x"CEE" => DATA <= x"20";
      when x"CEF" => DATA <= x"EB";
      when x"CF0" => DATA <= x"D0";
      when x"CF1" => DATA <= x"20";
      when x"CF2" => DATA <= x"24";
      when x"CF3" => DATA <= x"DD";
      when x"CF4" => DATA <= x"46";
      when x"CF5" => DATA <= x"6E";
      when x"CF6" => DATA <= x"90";
      when x"CF7" => DATA <= x"03";
      when x"CF8" => DATA <= x"20";
      when x"CF9" => DATA <= x"86";
      when x"CFA" => DATA <= x"DC";
      when x"CFB" => DATA <= x"46";
      when x"CFC" => DATA <= x"6E";
      when x"CFD" => DATA <= x"90";
      when x"CFE" => DATA <= x"06";
      when x"CFF" => DATA <= x"20";
      when x"D00" => DATA <= x"05";
      when x"D01" => DATA <= x"DD";
      when x"D02" => DATA <= x"4C";
      when x"D03" => DATA <= x"BF";
      when x"D04" => DATA <= x"D1";
      when x"D05" => DATA <= x"20";
      when x"D06" => DATA <= x"2C";
      when x"D07" => DATA <= x"D8";
      when x"D08" => DATA <= x"20";
      when x"D09" => DATA <= x"93";
      when x"D0A" => DATA <= x"DD";
      when x"D0B" => DATA <= x"20";
      when x"D0C" => DATA <= x"04";
      when x"D0D" => DATA <= x"D8";
      when x"D0E" => DATA <= x"C6";
      when x"D0F" => DATA <= x"61";
      when x"D10" => DATA <= x"A9";
      when x"D11" => DATA <= x"80";
      when x"D12" => DATA <= x"85";
      when x"D13" => DATA <= x"5F";
      when x"D14" => DATA <= x"20";
      when x"D15" => DATA <= x"41";
      when x"D16" => DATA <= x"D9";
      when x"D17" => DATA <= x"A9";
      when x"D18" => DATA <= x"A6";
      when x"D19" => DATA <= x"A0";
      when x"D1A" => DATA <= x"DD";
      when x"D1B" => DATA <= x"20";
      when x"D1C" => DATA <= x"27";
      when x"D1D" => DATA <= x"DC";
      when x"D1E" => DATA <= x"20";
      when x"D1F" => DATA <= x"A6";
      when x"D20" => DATA <= x"DB";
      when x"D21" => DATA <= x"4C";
      when x"D22" => DATA <= x"45";
      when x"D23" => DATA <= x"DA";
      when x"D24" => DATA <= x"A5";
      when x"D25" => DATA <= x"59";
      when x"D26" => DATA <= x"C9";
      when x"D27" => DATA <= x"98";
      when x"D28" => DATA <= x"B0";
      when x"D29" => DATA <= x"54";
      when x"D2A" => DATA <= x"20";
      when x"D2B" => DATA <= x"31";
      when x"D2C" => DATA <= x"D8";
      when x"D2D" => DATA <= x"20";
      when x"D2E" => DATA <= x"93";
      when x"D2F" => DATA <= x"DD";
      when x"D30" => DATA <= x"20";
      when x"D31" => DATA <= x"DC";
      when x"D32" => DATA <= x"DA";
      when x"D33" => DATA <= x"20";
      when x"D34" => DATA <= x"9A";
      when x"D35" => DATA <= x"D8";
      when x"D36" => DATA <= x"A5";
      when x"D37" => DATA <= x"5D";
      when x"D38" => DATA <= x"85";
      when x"D39" => DATA <= x"6E";
      when x"D3A" => DATA <= x"05";
      when x"D3B" => DATA <= x"5C";
      when x"D3C" => DATA <= x"05";
      when x"D3D" => DATA <= x"5B";
      when x"D3E" => DATA <= x"05";
      when x"D3F" => DATA <= x"5A";
      when x"D40" => DATA <= x"F0";
      when x"D41" => DATA <= x"3E";
      when x"D42" => DATA <= x"20";
      when x"D43" => DATA <= x"AC";
      when x"D44" => DATA <= x"D2";
      when x"D45" => DATA <= x"20";
      when x"D46" => DATA <= x"27";
      when x"D47" => DATA <= x"D8";
      when x"D48" => DATA <= x"20";
      when x"D49" => DATA <= x"86";
      when x"D4A" => DATA <= x"DD";
      when x"D4B" => DATA <= x"20";
      when x"D4C" => DATA <= x"45";
      when x"D4D" => DATA <= x"DA";
      when x"D4E" => DATA <= x"20";
      when x"D4F" => DATA <= x"AA";
      when x"D50" => DATA <= x"DB";
      when x"D51" => DATA <= x"20";
      when x"D52" => DATA <= x"3C";
      when x"D53" => DATA <= x"D9";
      when x"D54" => DATA <= x"20";
      when x"D55" => DATA <= x"3D";
      when x"D56" => DATA <= x"D8";
      when x"D57" => DATA <= x"20";
      when x"D58" => DATA <= x"A2";
      when x"D59" => DATA <= x"DB";
      when x"D5A" => DATA <= x"20";
      when x"D5B" => DATA <= x"E5";
      when x"D5C" => DATA <= x"D1";
      when x"D5D" => DATA <= x"20";
      when x"D5E" => DATA <= x"8A";
      when x"D5F" => DATA <= x"DD";
      when x"D60" => DATA <= x"20";
      when x"D61" => DATA <= x"45";
      when x"D62" => DATA <= x"DA";
      when x"D63" => DATA <= x"20";
      when x"D64" => DATA <= x"AA";
      when x"D65" => DATA <= x"DB";
      when x"D66" => DATA <= x"20";
      when x"D67" => DATA <= x"3C";
      when x"D68" => DATA <= x"D9";
      when x"D69" => DATA <= x"A5";
      when x"D6A" => DATA <= x"57";
      when x"D6B" => DATA <= x"10";
      when x"D6C" => DATA <= x"12";
      when x"D6D" => DATA <= x"20";
      when x"D6E" => DATA <= x"8A";
      when x"D6F" => DATA <= x"DD";
      when x"D70" => DATA <= x"20";
      when x"D71" => DATA <= x"33";
      when x"D72" => DATA <= x"D9";
      when x"D73" => DATA <= x"20";
      when x"D74" => DATA <= x"86";
      when x"D75" => DATA <= x"DD";
      when x"D76" => DATA <= x"20";
      when x"D77" => DATA <= x"33";
      when x"D78" => DATA <= x"D9";
      when x"D79" => DATA <= x"C6";
      when x"D7A" => DATA <= x"6E";
      when x"D7B" => DATA <= x"4C";
      when x"D7C" => DATA <= x"69";
      when x"D7D" => DATA <= x"DD";
      when x"D7E" => DATA <= x"00";
      when x"D7F" => DATA <= x"60";
      when x"D80" => DATA <= x"20";
      when x"D81" => DATA <= x"DA";
      when x"D82" => DATA <= x"D2";
      when x"D83" => DATA <= x"4C";
      when x"D84" => DATA <= x"69";
      when x"D85" => DATA <= x"DD";
      when x"D86" => DATA <= x"A9";
      when x"D87" => DATA <= x"97";
      when x"D88" => DATA <= x"D0";
      when x"D89" => DATA <= x"02";
      when x"D8A" => DATA <= x"A9";
      when x"D8B" => DATA <= x"9C";
      when x"D8C" => DATA <= x"85";
      when x"D8D" => DATA <= x"6F";
      when x"D8E" => DATA <= x"A9";
      when x"D8F" => DATA <= x"DD";
      when x"D90" => DATA <= x"85";
      when x"D91" => DATA <= x"70";
      when x"D92" => DATA <= x"60";
      when x"D93" => DATA <= x"A9";
      when x"D94" => DATA <= x"A1";
      when x"D95" => DATA <= x"D0";
      when x"D96" => DATA <= x"F5";
      when x"D97" => DATA <= x"81";
      when x"D98" => DATA <= x"C9";
      when x"D99" => DATA <= x"00";
      when x"D9A" => DATA <= x"00";
      when x"D9B" => DATA <= x"00";
      when x"D9C" => DATA <= x"75";
      when x"D9D" => DATA <= x"FD";
      when x"D9E" => DATA <= x"AA";
      when x"D9F" => DATA <= x"22";
      when x"DA0" => DATA <= x"17";
      when x"DA1" => DATA <= x"81";
      when x"DA2" => DATA <= x"49";
      when x"DA3" => DATA <= x"0F";
      when x"DA4" => DATA <= x"DA";
      when x"DA5" => DATA <= x"A2";
      when x"DA6" => DATA <= x"08";
      when x"DA7" => DATA <= x"84";
      when x"DA8" => DATA <= x"04";
      when x"DA9" => DATA <= x"C7";
      when x"DAA" => DATA <= x"3C";
      when x"DAB" => DATA <= x"FB";
      when x"DAC" => DATA <= x"81";
      when x"DAD" => DATA <= x"E0";
      when x"DAE" => DATA <= x"4F";
      when x"DAF" => DATA <= x"5D";
      when x"DB0" => DATA <= x"AD";
      when x"DB1" => DATA <= x"82";
      when x"DB2" => DATA <= x"80";
      when x"DB3" => DATA <= x"00";
      when x"DB4" => DATA <= x"69";
      when x"DB5" => DATA <= x"B8";
      when x"DB6" => DATA <= x"82";
      when x"DB7" => DATA <= x"5B";
      when x"DB8" => DATA <= x"CF";
      when x"DB9" => DATA <= x"1D";
      when x"DBA" => DATA <= x"B5";
      when x"DBB" => DATA <= x"82";
      when x"DBC" => DATA <= x"BF";
      when x"DBD" => DATA <= x"CE";
      when x"DBE" => DATA <= x"82";
      when x"DBF" => DATA <= x"1E";
      when x"DC0" => DATA <= x"82";
      when x"DC1" => DATA <= x"45";
      when x"DC2" => DATA <= x"44";
      when x"DC3" => DATA <= x"7F";
      when x"DC4" => DATA <= x"32";
      when x"DC5" => DATA <= x"7F";
      when x"DC6" => DATA <= x"62";
      when x"DC7" => DATA <= x"44";
      when x"DC8" => DATA <= x"5A";
      when x"DC9" => DATA <= x"D2";
      when x"DCA" => DATA <= x"83";
      when x"DCB" => DATA <= x"82";
      when x"DCC" => DATA <= x"14";
      when x"DCD" => DATA <= x"8A";
      when x"DCE" => DATA <= x"27";
      when x"DCF" => DATA <= x"80";
      when x"DD0" => DATA <= x"66";
      when x"DD1" => DATA <= x"7B";
      when x"DD2" => DATA <= x"21";
      when x"DD3" => DATA <= x"4D";
      when x"DD4" => DATA <= x"20";
      when x"DD5" => DATA <= x"EB";
      when x"DD6" => DATA <= x"D0";
      when x"DD7" => DATA <= x"A5";
      when x"DD8" => DATA <= x"59";
      when x"DD9" => DATA <= x"C9";
      when x"DDA" => DATA <= x"87";
      when x"DDB" => DATA <= x"90";
      when x"DDC" => DATA <= x"10";
      when x"DDD" => DATA <= x"D0";
      when x"DDE" => DATA <= x"06";
      when x"DDF" => DATA <= x"A5";
      when x"DE0" => DATA <= x"5A";
      when x"DE1" => DATA <= x"C9";
      when x"DE2" => DATA <= x"B3";
      when x"DE3" => DATA <= x"90";
      when x"DE4" => DATA <= x"08";
      when x"DE5" => DATA <= x"A5";
      when x"DE6" => DATA <= x"57";
      when x"DE7" => DATA <= x"10";
      when x"DE8" => DATA <= x"03";
      when x"DE9" => DATA <= x"4C";
      when x"DEA" => DATA <= x"A4";
      when x"DEB" => DATA <= x"DA";
      when x"DEC" => DATA <= x"00";
      when x"DED" => DATA <= x"A5";
      when x"DEE" => DATA <= x"59";
      when x"DEF" => DATA <= x"C9";
      when x"DF0" => DATA <= x"80";
      when x"DF1" => DATA <= x"90";
      when x"DF2" => DATA <= x"29";
      when x"DF3" => DATA <= x"20";
      when x"DF4" => DATA <= x"9A";
      when x"DF5" => DATA <= x"D8";
      when x"DF6" => DATA <= x"20";
      when x"DF7" => DATA <= x"E2";
      when x"DF8" => DATA <= x"D8";
      when x"DF9" => DATA <= x"A5";
      when x"DFA" => DATA <= x"5D";
      when x"DFB" => DATA <= x"85";
      when x"DFC" => DATA <= x"6E";
      when x"DFD" => DATA <= x"20";
      when x"DFE" => DATA <= x"13";
      when x"DFF" => DATA <= x"D9";
      when x"E00" => DATA <= x"20";
      when x"E01" => DATA <= x"1C";
      when x"E02" => DATA <= x"DE";
      when x"E03" => DATA <= x"20";
      when x"E04" => DATA <= x"2C";
      when x"E05" => DATA <= x"D8";
      when x"E06" => DATA <= x"A9";
      when x"E07" => DATA <= x"23";
      when x"E08" => DATA <= x"85";
      when x"E09" => DATA <= x"6F";
      when x"E0A" => DATA <= x"A9";
      when x"E0B" => DATA <= x"DE";
      when x"E0C" => DATA <= x"85";
      when x"E0D" => DATA <= x"70";
      when x"E0E" => DATA <= x"20";
      when x"E0F" => DATA <= x"E5";
      when x"E10" => DATA <= x"D1";
      when x"E11" => DATA <= x"A5";
      when x"E12" => DATA <= x"6E";
      when x"E13" => DATA <= x"20";
      when x"E14" => DATA <= x"51";
      when x"E15" => DATA <= x"DE";
      when x"E16" => DATA <= x"20";
      when x"E17" => DATA <= x"A6";
      when x"E18" => DATA <= x"DB";
      when x"E19" => DATA <= x"4C";
      when x"E1A" => DATA <= x"45";
      when x"E1B" => DATA <= x"DA";
      when x"E1C" => DATA <= x"A9";
      when x"E1D" => DATA <= x"28";
      when x"E1E" => DATA <= x"A0";
      when x"E1F" => DATA <= x"DE";
      when x"E20" => DATA <= x"4C";
      when x"E21" => DATA <= x"27";
      when x"E22" => DATA <= x"DC";
      when x"E23" => DATA <= x"82";
      when x"E24" => DATA <= x"2D";
      when x"E25" => DATA <= x"F8";
      when x"E26" => DATA <= x"54";
      when x"E27" => DATA <= x"58";
      when x"E28" => DATA <= x"07";
      when x"E29" => DATA <= x"83";
      when x"E2A" => DATA <= x"E0";
      when x"E2B" => DATA <= x"20";
      when x"E2C" => DATA <= x"86";
      when x"E2D" => DATA <= x"5B";
      when x"E2E" => DATA <= x"82";
      when x"E2F" => DATA <= x"80";
      when x"E30" => DATA <= x"53";
      when x"E31" => DATA <= x"93";
      when x"E32" => DATA <= x"B8";
      when x"E33" => DATA <= x"83";
      when x"E34" => DATA <= x"20";
      when x"E35" => DATA <= x"00";
      when x"E36" => DATA <= x"06";
      when x"E37" => DATA <= x"A1";
      when x"E38" => DATA <= x"82";
      when x"E39" => DATA <= x"00";
      when x"E3A" => DATA <= x"00";
      when x"E3B" => DATA <= x"21";
      when x"E3C" => DATA <= x"63";
      when x"E3D" => DATA <= x"82";
      when x"E3E" => DATA <= x"C0";
      when x"E3F" => DATA <= x"00";
      when x"E40" => DATA <= x"00";
      when x"E41" => DATA <= x"02";
      when x"E42" => DATA <= x"82";
      when x"E43" => DATA <= x"80";
      when x"E44" => DATA <= x"00";
      when x"E45" => DATA <= x"00";
      when x"E46" => DATA <= x"0C";
      when x"E47" => DATA <= x"81";
      when x"E48" => DATA <= x"00";
      when x"E49" => DATA <= x"00";
      when x"E4A" => DATA <= x"00";
      when x"E4B" => DATA <= x"00";
      when x"E4C" => DATA <= x"81";
      when x"E4D" => DATA <= x"00";
      when x"E4E" => DATA <= x"00";
      when x"E4F" => DATA <= x"00";
      when x"E50" => DATA <= x"00";
      when x"E51" => DATA <= x"AA";
      when x"E52" => DATA <= x"10";
      when x"E53" => DATA <= x"09";
      when x"E54" => DATA <= x"CA";
      when x"E55" => DATA <= x"8A";
      when x"E56" => DATA <= x"49";
      when x"E57" => DATA <= x"FF";
      when x"E58" => DATA <= x"48";
      when x"E59" => DATA <= x"20";
      when x"E5A" => DATA <= x"AE";
      when x"E5B" => DATA <= x"DA";
      when x"E5C" => DATA <= x"68";
      when x"E5D" => DATA <= x"48";
      when x"E5E" => DATA <= x"20";
      when x"E5F" => DATA <= x"31";
      when x"E60" => DATA <= x"D8";
      when x"E61" => DATA <= x"20";
      when x"E62" => DATA <= x"8D";
      when x"E63" => DATA <= x"DE";
      when x"E64" => DATA <= x"68";
      when x"E65" => DATA <= x"F0";
      when x"E66" => DATA <= x"0A";
      when x"E67" => DATA <= x"38";
      when x"E68" => DATA <= x"E9";
      when x"E69" => DATA <= x"01";
      when x"E6A" => DATA <= x"48";
      when x"E6B" => DATA <= x"20";
      when x"E6C" => DATA <= x"45";
      when x"E6D" => DATA <= x"DA";
      when x"E6E" => DATA <= x"4C";
      when x"E6F" => DATA <= x"64";
      when x"E70" => DATA <= x"DE";
      when x"E71" => DATA <= x"60";
      when x"E72" => DATA <= x"20";
      when x"E73" => DATA <= x"EB";
      when x"E74" => DATA <= x"D0";
      when x"E75" => DATA <= x"A5";
      when x"E76" => DATA <= x"57";
      when x"E77" => DATA <= x"10";
      when x"E78" => DATA <= x"0A";
      when x"E79" => DATA <= x"A9";
      when x"E7A" => DATA <= x"00";
      when x"E7B" => DATA <= x"85";
      when x"E7C" => DATA <= x"57";
      when x"E7D" => DATA <= x"20";
      when x"E7E" => DATA <= x"83";
      when x"E7F" => DATA <= x"DE";
      when x"E80" => DATA <= x"4C";
      when x"E81" => DATA <= x"BF";
      when x"E82" => DATA <= x"D1";
      when x"E83" => DATA <= x"A5";
      when x"E84" => DATA <= x"59";
      when x"E85" => DATA <= x"C9";
      when x"E86" => DATA <= x"81";
      when x"E87" => DATA <= x"90";
      when x"E88" => DATA <= x"33";
      when x"E89" => DATA <= x"C9";
      when x"E8A" => DATA <= x"85";
      when x"E8B" => DATA <= x"90";
      when x"E8C" => DATA <= x"0B";
      when x"E8D" => DATA <= x"20";
      when x"E8E" => DATA <= x"A4";
      when x"E8F" => DATA <= x"DA";
      when x"E90" => DATA <= x"A0";
      when x"E91" => DATA <= x"80";
      when x"E92" => DATA <= x"84";
      when x"E93" => DATA <= x"5A";
      when x"E94" => DATA <= x"C8";
      when x"E95" => DATA <= x"84";
      when x"E96" => DATA <= x"59";
      when x"E97" => DATA <= x"60";
      when x"E98" => DATA <= x"E6";
      when x"E99" => DATA <= x"59";
      when x"E9A" => DATA <= x"A9";
      when x"E9B" => DATA <= x"80";
      when x"E9C" => DATA <= x"85";
      when x"E9D" => DATA <= x"57";
      when x"E9E" => DATA <= x"20";
      when x"E9F" => DATA <= x"D7";
      when x"EA0" => DATA <= x"DD";
      when x"EA1" => DATA <= x"20";
      when x"EA2" => DATA <= x"31";
      when x"EA3" => DATA <= x"D8";
      when x"EA4" => DATA <= x"20";
      when x"EA5" => DATA <= x"8D";
      when x"EA6" => DATA <= x"DE";
      when x"EA7" => DATA <= x"20";
      when x"EA8" => DATA <= x"3C";
      when x"EA9" => DATA <= x"D9";
      when x"EAA" => DATA <= x"20";
      when x"EAB" => DATA <= x"27";
      when x"EAC" => DATA <= x"D8";
      when x"EAD" => DATA <= x"20";
      when x"EAE" => DATA <= x"8D";
      when x"EAF" => DATA <= x"DE";
      when x"EB0" => DATA <= x"20";
      when x"EB1" => DATA <= x"AA";
      when x"EB2" => DATA <= x"DB";
      when x"EB3" => DATA <= x"20";
      when x"EB4" => DATA <= x"33";
      when x"EB5" => DATA <= x"D9";
      when x"EB6" => DATA <= x"20";
      when x"EB7" => DATA <= x"A2";
      when x"EB8" => DATA <= x"DB";
      when x"EB9" => DATA <= x"4C";
      when x"EBA" => DATA <= x"DC";
      when x"EBB" => DATA <= x"DA";
      when x"EBC" => DATA <= x"20";
      when x"EBD" => DATA <= x"2C";
      when x"EBE" => DATA <= x"D8";
      when x"EBF" => DATA <= x"20";
      when x"EC0" => DATA <= x"8D";
      when x"EC1" => DATA <= x"DE";
      when x"EC2" => DATA <= x"C6";
      when x"EC3" => DATA <= x"59";
      when x"EC4" => DATA <= x"20";
      when x"EC5" => DATA <= x"33";
      when x"EC6" => DATA <= x"D9";
      when x"EC7" => DATA <= x"A9";
      when x"EC8" => DATA <= x"D4";
      when x"EC9" => DATA <= x"A0";
      when x"ECA" => DATA <= x"DE";
      when x"ECB" => DATA <= x"20";
      when x"ECC" => DATA <= x"27";
      when x"ECD" => DATA <= x"DC";
      when x"ECE" => DATA <= x"20";
      when x"ECF" => DATA <= x"A6";
      when x"ED0" => DATA <= x"DB";
      when x"ED1" => DATA <= x"4C";
      when x"ED2" => DATA <= x"45";
      when x"ED3" => DATA <= x"DA";
      when x"ED4" => DATA <= x"08";
      when x"ED5" => DATA <= x"7E";
      when x"ED6" => DATA <= x"85";
      when x"ED7" => DATA <= x"51";
      when x"ED8" => DATA <= x"B3";
      when x"ED9" => DATA <= x"0C";
      when x"EDA" => DATA <= x"86";
      when x"EDB" => DATA <= x"DE";
      when x"EDC" => DATA <= x"B0";
      when x"EDD" => DATA <= x"7D";
      when x"EDE" => DATA <= x"73";
      when x"EDF" => DATA <= x"7C";
      when x"EE0" => DATA <= x"23";
      when x"EE1" => DATA <= x"D8";
      when x"EE2" => DATA <= x"E9";
      when x"EE3" => DATA <= x"9A";
      when x"EE4" => DATA <= x"87";
      when x"EE5" => DATA <= x"34";
      when x"EE6" => DATA <= x"82";
      when x"EE7" => DATA <= x"1D";
      when x"EE8" => DATA <= x"80";
      when x"EE9" => DATA <= x"81";
      when x"EEA" => DATA <= x"9A";
      when x"EEB" => DATA <= x"20";
      when x"EEC" => DATA <= x"6C";
      when x"EED" => DATA <= x"ED";
      when x"EEE" => DATA <= x"81";
      when x"EEF" => DATA <= x"BD";
      when x"EF0" => DATA <= x"32";
      when x"EF1" => DATA <= x"34";
      when x"EF2" => DATA <= x"2E";
      when x"EF3" => DATA <= x"7F";
      when x"EF4" => DATA <= x"5D";
      when x"EF5" => DATA <= x"46";
      when x"EF6" => DATA <= x"87";
      when x"EF7" => DATA <= x"B4";
      when x"EF8" => DATA <= x"82";
      when x"EF9" => DATA <= x"68";
      when x"EFA" => DATA <= x"3E";
      when x"EFB" => DATA <= x"43";
      when x"EFC" => DATA <= x"F7";
      when x"EFD" => DATA <= x"80";
      when x"EFE" => DATA <= x"6C";
      when x"EFF" => DATA <= x"9A";
      when x"F00" => DATA <= x"9E";
      when x"F01" => DATA <= x"BB";
      when x"F02" => DATA <= x"20";
      when x"F03" => DATA <= x"C8";
      when x"F04" => DATA <= x"C3";
      when x"F05" => DATA <= x"A5";
      when x"F06" => DATA <= x"52";
      when x"F07" => DATA <= x"29";
      when x"F08" => DATA <= x"03";
      when x"F09" => DATA <= x"A8";
      when x"F0A" => DATA <= x"B9";
      when x"F0B" => DATA <= x"4E";
      when x"F0C" => DATA <= x"DF";
      when x"F0D" => DATA <= x"8D";
      when x"F0E" => DATA <= x"FD";
      when x"F0F" => DATA <= x"03";
      when x"F10" => DATA <= x"AD";
      when x"F11" => DATA <= x"00";
      when x"F12" => DATA <= x"B0";
      when x"F13" => DATA <= x"29";
      when x"F14" => DATA <= x"F0";
      when x"F15" => DATA <= x"C9";
      when x"F16" => DATA <= x"70";
      when x"F17" => DATA <= x"D0";
      when x"F18" => DATA <= x"0C";
      when x"F19" => DATA <= x"A9";
      when x"F1A" => DATA <= x"00";
      when x"F1B" => DATA <= x"A8";
      when x"F1C" => DATA <= x"99";
      when x"F1D" => DATA <= x"00";
      when x"F1E" => DATA <= x"86";
      when x"F1F" => DATA <= x"99";
      when x"F20" => DATA <= x"00";
      when x"F21" => DATA <= x"87";
      when x"F22" => DATA <= x"88";
      when x"F23" => DATA <= x"D0";
      when x"F24" => DATA <= x"F7";
      when x"F25" => DATA <= x"AD";
      when x"F26" => DATA <= x"00";
      when x"F27" => DATA <= x"B0";
      when x"F28" => DATA <= x"29";
      when x"F29" => DATA <= x"DF";
      when x"F2A" => DATA <= x"8D";
      when x"F2B" => DATA <= x"00";
      when x"F2C" => DATA <= x"B0";
      when x"F2D" => DATA <= x"2A";
      when x"F2E" => DATA <= x"2A";
      when x"F2F" => DATA <= x"2A";
      when x"F30" => DATA <= x"29";
      when x"F31" => DATA <= x"03";
      when x"F32" => DATA <= x"A8";
      when x"F33" => DATA <= x"B9";
      when x"F34" => DATA <= x"42";
      when x"F35" => DATA <= x"DF";
      when x"F36" => DATA <= x"8D";
      when x"F37" => DATA <= x"FE";
      when x"F38" => DATA <= x"03";
      when x"F39" => DATA <= x"B9";
      when x"F3A" => DATA <= x"46";
      when x"F3B" => DATA <= x"DF";
      when x"F3C" => DATA <= x"8D";
      when x"F3D" => DATA <= x"FF";
      when x"F3E" => DATA <= x"03";
      when x"F3F" => DATA <= x"4C";
      when x"F40" => DATA <= x"58";
      when x"F41" => DATA <= x"C5";
      when x"F42" => DATA <= x"52";
      when x"F43" => DATA <= x"70";
      when x"F44" => DATA <= x"88";
      when x"F45" => DATA <= x"A0";
      when x"F46" => DATA <= x"DF";
      when x"F47" => DATA <= x"DF";
      when x"F48" => DATA <= x"DF";
      when x"F49" => DATA <= x"DF";
      when x"F4A" => DATA <= x"3F";
      when x"F4B" => DATA <= x"CF";
      when x"F4C" => DATA <= x"F3";
      when x"F4D" => DATA <= x"FC";
      when x"F4E" => DATA <= x"00";
      when x"F4F" => DATA <= x"55";
      when x"F50" => DATA <= x"AA";
      when x"F51" => DATA <= x"FF";
      when x"F52" => DATA <= x"A5";
      when x"F53" => DATA <= x"5B";
      when x"F54" => DATA <= x"05";
      when x"F55" => DATA <= x"5D";
      when x"F56" => DATA <= x"D0";
      when x"F57" => DATA <= x"47";
      when x"F58" => DATA <= x"A5";
      when x"F59" => DATA <= x"5A";
      when x"F5A" => DATA <= x"C9";
      when x"F5B" => DATA <= x"40";
      when x"F5C" => DATA <= x"B0";
      when x"F5D" => DATA <= x"41";
      when x"F5E" => DATA <= x"4A";
      when x"F5F" => DATA <= x"4A";
      when x"F60" => DATA <= x"85";
      when x"F61" => DATA <= x"5F";
      when x"F62" => DATA <= x"A0";
      when x"F63" => DATA <= x"00";
      when x"F64" => DATA <= x"84";
      when x"F65" => DATA <= x"60";
      when x"F66" => DATA <= x"A9";
      when x"F67" => DATA <= x"3F";
      when x"F68" => DATA <= x"38";
      when x"F69" => DATA <= x"E5";
      when x"F6A" => DATA <= x"5C";
      when x"F6B" => DATA <= x"C9";
      when x"F6C" => DATA <= x"40";
      when x"F6D" => DATA <= x"90";
      when x"F6E" => DATA <= x"4F";
      when x"F6F" => DATA <= x"60";
      when x"F70" => DATA <= x"A5";
      when x"F71" => DATA <= x"5B";
      when x"F72" => DATA <= x"05";
      when x"F73" => DATA <= x"5D";
      when x"F74" => DATA <= x"D0";
      when x"F75" => DATA <= x"29";
      when x"F76" => DATA <= x"A5";
      when x"F77" => DATA <= x"5A";
      when x"F78" => DATA <= x"30";
      when x"F79" => DATA <= x"25";
      when x"F7A" => DATA <= x"4A";
      when x"F7B" => DATA <= x"4A";
      when x"F7C" => DATA <= x"85";
      when x"F7D" => DATA <= x"5F";
      when x"F7E" => DATA <= x"A9";
      when x"F7F" => DATA <= x"3F";
      when x"F80" => DATA <= x"38";
      when x"F81" => DATA <= x"E5";
      when x"F82" => DATA <= x"5C";
      when x"F83" => DATA <= x"C9";
      when x"F84" => DATA <= x"40";
      when x"F85" => DATA <= x"90";
      when x"F86" => DATA <= x"30";
      when x"F87" => DATA <= x"60";
      when x"F88" => DATA <= x"A5";
      when x"F89" => DATA <= x"5B";
      when x"F8A" => DATA <= x"05";
      when x"F8B" => DATA <= x"5D";
      when x"F8C" => DATA <= x"D0";
      when x"F8D" => DATA <= x"11";
      when x"F8E" => DATA <= x"A5";
      when x"F8F" => DATA <= x"5A";
      when x"F90" => DATA <= x"30";
      when x"F91" => DATA <= x"0D";
      when x"F92" => DATA <= x"4A";
      when x"F93" => DATA <= x"4A";
      when x"F94" => DATA <= x"85";
      when x"F95" => DATA <= x"5F";
      when x"F96" => DATA <= x"A9";
      when x"F97" => DATA <= x"5F";
      when x"F98" => DATA <= x"38";
      when x"F99" => DATA <= x"E5";
      when x"F9A" => DATA <= x"5C";
      when x"F9B" => DATA <= x"C9";
      when x"F9C" => DATA <= x"60";
      when x"F9D" => DATA <= x"90";
      when x"F9E" => DATA <= x"18";
      when x"F9F" => DATA <= x"60";
      when x"FA0" => DATA <= x"A5";
      when x"FA1" => DATA <= x"5B";
      when x"FA2" => DATA <= x"05";
      when x"FA3" => DATA <= x"5D";
      when x"FA4" => DATA <= x"D0";
      when x"FA5" => DATA <= x"F9";
      when x"FA6" => DATA <= x"A5";
      when x"FA7" => DATA <= x"5A";
      when x"FA8" => DATA <= x"30";
      when x"FA9" => DATA <= x"F5";
      when x"FAA" => DATA <= x"4A";
      when x"FAB" => DATA <= x"4A";
      when x"FAC" => DATA <= x"85";
      when x"FAD" => DATA <= x"5F";
      when x"FAE" => DATA <= x"A9";
      when x"FAF" => DATA <= x"BF";
      when x"FB0" => DATA <= x"38";
      when x"FB1" => DATA <= x"E5";
      when x"FB2" => DATA <= x"5C";
      when x"FB3" => DATA <= x"C9";
      when x"FB4" => DATA <= x"C0";
      when x"FB5" => DATA <= x"B0";
      when x"FB6" => DATA <= x"E8";
      when x"FB7" => DATA <= x"A0";
      when x"FB8" => DATA <= x"00";
      when x"FB9" => DATA <= x"84";
      when x"FBA" => DATA <= x"60";
      when x"FBB" => DATA <= x"0A";
      when x"FBC" => DATA <= x"26";
      when x"FBD" => DATA <= x"60";
      when x"FBE" => DATA <= x"0A";
      when x"FBF" => DATA <= x"26";
      when x"FC0" => DATA <= x"60";
      when x"FC1" => DATA <= x"0A";
      when x"FC2" => DATA <= x"26";
      when x"FC3" => DATA <= x"60";
      when x"FC4" => DATA <= x"0A";
      when x"FC5" => DATA <= x"26";
      when x"FC6" => DATA <= x"60";
      when x"FC7" => DATA <= x"0A";
      when x"FC8" => DATA <= x"26";
      when x"FC9" => DATA <= x"60";
      when x"FCA" => DATA <= x"65";
      when x"FCB" => DATA <= x"5F";
      when x"FCC" => DATA <= x"85";
      when x"FCD" => DATA <= x"5F";
      when x"FCE" => DATA <= x"A5";
      when x"FCF" => DATA <= x"60";
      when x"FD0" => DATA <= x"69";
      when x"FD1" => DATA <= x"80";
      when x"FD2" => DATA <= x"85";
      when x"FD3" => DATA <= x"60";
      when x"FD4" => DATA <= x"A5";
      when x"FD5" => DATA <= x"5A";
      when x"FD6" => DATA <= x"29";
      when x"FD7" => DATA <= x"03";
      when x"FD8" => DATA <= x"AA";
      when x"FD9" => DATA <= x"BD";
      when x"FDA" => DATA <= x"4A";
      when x"FDB" => DATA <= x"DF";
      when x"FDC" => DATA <= x"A6";
      when x"FDD" => DATA <= x"5E";
      when x"FDE" => DATA <= x"CA";
      when x"FDF" => DATA <= x"F0";
      when x"FE0" => DATA <= x"0F";
      when x"FE1" => DATA <= x"CA";
      when x"FE2" => DATA <= x"F0";
      when x"FE3" => DATA <= x"05";
      when x"FE4" => DATA <= x"31";
      when x"FE5" => DATA <= x"5F";
      when x"FE6" => DATA <= x"91";
      when x"FE7" => DATA <= x"5F";
      when x"FE8" => DATA <= x"60";
      when x"FE9" => DATA <= x"49";
      when x"FEA" => DATA <= x"FF";
      when x"FEB" => DATA <= x"51";
      when x"FEC" => DATA <= x"5F";
      when x"FED" => DATA <= x"91";
      when x"FEE" => DATA <= x"5F";
      when x"FEF" => DATA <= x"60";
      when x"FF0" => DATA <= x"AA";
      when x"FF1" => DATA <= x"31";
      when x"FF2" => DATA <= x"5F";
      when x"FF3" => DATA <= x"91";
      when x"FF4" => DATA <= x"5F";
      when x"FF5" => DATA <= x"8A";
      when x"FF6" => DATA <= x"49";
      when x"FF7" => DATA <= x"FF";
      when x"FF8" => DATA <= x"2D";
      when x"FF9" => DATA <= x"FD";
      when x"FFA" => DATA <= x"03";
      when x"FFB" => DATA <= x"11";
      when x"FFC" => DATA <= x"5F";
      when x"FFD" => DATA <= x"91";
      when x"FFE" => DATA <= x"5F";
      when x"FFF" => DATA <= x"60";
      when others => DATA <= (others => '0');
    end case;
  end process;
end RTL;
